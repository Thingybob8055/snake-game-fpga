library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity snake is
    Port ( clk_100mhz : in STD_LOGIC;					--  master clock 100MHz
		   pixel_clk : in STD_LOGIC;					-- pixel clock
		   update : in STD_LOGIC;						-- signal to update the food position
		   clk_500hz : in STD_LOGIC;					-- 500Hz clock
		   xCount : in unsigned(10 downto 0);			-- x position from horizontal counter of vga driver
		   yCount : in unsigned(10 downto 0);			-- y position from vertical counter of vga driver
		   rand_X : in unsigned(6 downto 0);			-- random x position for the food
		   rand_Y : in unsigned(6 downto 0);			-- random y position for the food
           switch : in STD_LOGIC_VECTOR(7 downto 0);	-- switches 0-7
           btn_up : in STD_LOGIC;						-- up button
           btn_left : in STD_LOGIC;						-- left button
           btn_right : in STD_LOGIC;					-- right button
           btn_down : in STD_LOGIC;						-- down button
		   display : in STD_LOGIC;						-- display signal to enable rgb when blanking is off
           led : out STD_LOGIC_VECTOR(7 downto 0);		-- leds 0-7
           vgared : out STD_LOGIC_VECTOR(3 downto 0);	-- vga red
           vgagreen : out STD_LOGIC_VECTOR(3 downto 0);	-- vga green
           vgablue : out STD_LOGIC_VECTOR(3 downto 0);	-- vga blue
		   seg  : out std_logic_vector (6 downto 0); 	-- 7-segment display
           dp   : out std_logic; 						-- 7-segment display decimal point
           an   : out std_logic_vector (3 downto 0)		-- 7-segment display anodes
         );
end snake;

architecture Behavioral of snake is
    constant SIZE_INCREMENT : integer := 4;   -- size increment for the snake body
    
    signal size : unsigned(6 downto 0);	    -- keep track of the size of the snake
    signal pearX : unsigned(6 downto 0) := "0101000"; 
    signal pearY : unsigned(6 downto 0) := "0001010";
    signal game_over : std_logic;  -- signal to indicate game over
    signal border : std_logic; -- signal to draw border and food

    type snake_array is array (0 to 127) of unsigned(6 downto 0);  -- array to keep track of the snake body
    -- type snakeY_array is array (0 to 127) of unsigned(6 downto 0);

    signal snakeX : snake_array;	-- snake x positions
    signal snakeY : snake_array;	-- snake y positions

    signal snakeBody : unsigned(127 downto 0);  -- vector to render the snake body
    signal direction : std_logic_vector(3 downto 0) := "0001";

    signal count : integer;  -- counter to keep track of the snake body in the for loops

    signal start : std_logic;  -- signal to start the game
    
	-- rick astley never gonna give you up GIF
    type color_gif_sprite is array (0 to 31, 0 to 47, 0 to 26) of std_logic_vector(0 to 11);
	constant COLOR_GIF_ROM : color_gif_sprite := (

		(	("100001111001","100001111001","100110001010","100001111001","100001111001","100010001010","100110011011","100110001010","100010001010","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100001111001","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100010001010","100010001010","100010001010","100010001010","100001111001","100001111001","100001111001","100010001010","100001111001","100001111001","100110001010","100110011011","100110011011","100110001010","100010001010","100010001010","100010001010","100010001010","100010001010","100010001010","100110001010","100110001010","100001111000","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100010001010","100010001010","100001111001","100001111001","100110011011","101010011011","101010101100","101010101100","101010011011","100110001010","100110001010","100110011011","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110011011","101010101100","101010011011","100110011011","100010001010","100010001010","100001111001","100110011011","101010011011","101010101100","101010101100","101010101100","101010101100","100110001010","100010001010","100010001010","100110001010","100110001010","100110011011","100010001010","100001111001","100001111001"),
		("101110101100","100110011011","100110001010","100110011011","100110011011","100110011011","101010101100","101010101100","100110011011","100110011011","100010001010","100110001010","101010011011","101010101100","101010101100","101010101100","101110101100","101110101100","101010011011","100110011011","100110001010","101010101100","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110001010","100110001010","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001010","100010001010","101010101100","101010101100","101010101100","101110101100","101110101100","101110101100","101010101100","100110011011","100110001010","101010011011","101010011011","100110001010","100010001010","100001111001","100001111001"),
		("100110001010","101010101100","100110011011","100110011011","100110011011","101010101100","100110001010","100010001010","100010001010","100010001010","100001111001","100010001010","100010001010","101010101100","101010101100","101110101100","101110101100","101010101100","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100110001010","100001111001"),
		("101010101100","101110101100","100110011011","100110011011","100110011011","100110011011","100110001010","101010101100","101110101100","101010101100","101010101100","100001111001","100010001010","101010011011","101010101100","101010101100","101010101100","101010011011","100110001010","100010001010","101010011011","101010011011","100010001010","100001111001","100001111001","100110001010","100001111001"),
		("101110101100","101110111101","100110011011","100110011011","100110011011","100110011011","101010011011","101110101100","101110101100","101010101100","101010101100","100110001010","100010001010","100010001010","100101100111","100001000011","100101100101","100101100111","100110001010","101010101100","101010101100","101010011011","101010011011","100010001010","100001111001","100001111001","100001111001"),
		("101110101100","101110111101","100110011011","100110011011","100110011011","101010101100","101110101100","101110101100","101010101100","101010101100","101010101100","100110001010","101010011010","100101100111","010100100010","010100100010","010100100010","011100110011","011000110011","101010011010","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("100110011011","101110101100","100110011011","100110011011","100110011011","100110011011","101110111101","101110111101","101110101100","101010011011","101010011011","100101111000","100101100101","100001000011","010100100010","010000100001","010000100001","010100100010","011000110011","011000110011","100110001001","100110011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","101110101100","101110101100","101110101100","101110101100","101010101100","101010011011","100101111000","100001000011","011100110011","010000100001","010000100010","010000100010","010000100001","010000100001","010000100001","011000110011","101010011010","100110011011","100110011011","100010001010","100001111001","100001111001"),
		("101110101100","100110011011","100110011011","100110011011","100110011011","101110101100","101110101100","101110101100","101110101100","101110101100","101010101100","100101100111","010100100010","011101000100","011101000100","100001010101","011000110011","010100100010","010100100010","010100100010","011000110011","101010011011","101010011011","100110011011","100110011011","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110011011","100110001010","100110011011","100110001010","101010101100","101010101100","101010011011","101010011010","100001000011","011000110100","100001000101","011101000101","100101100110","100101100110","100101100111","100101100111","011000110011","011000110100","101010011011","101010011011","100110011011","100110011011","100001111001","100001111001"),
		("101110101100","101110101100","100110001010","100110001010","100110011011","100110001010","100110001010","101010101100","101010101100","101010011011","100101111000","011100110011","011101000100","011100110011","011101000100","100101100110","100101100110","100101100110","100001010110","011101000101","100101111000","101010011011","101010011011","101010011010","100001111001","100001111001","100001111001"),
		("101110101100","101010101100","100110001010","100110001010","101010011011","101010101100","100110001010","100110001010","100010001010","100010001010","100001000101","100101100101","100001010101","011000110100","011000110100","011101000100","100001010110","100101100110","100001010110","011101000100","100110001001","101010101100","101010011011","100001111001","100001111001","100110001010","100001111001"),
		("101110101100","101010101100","100110001010","100110001010","100110011011","100110001010","100010001010","100010001010","100010001010","100001111001","100001000101","100101100101","100001010101","100001010110","100001010110","100001010101","100001010110","011000110100","100001010101","100001010110","100110001001","100010001010","100010001010","100001111001","100001111001","100110001010","100001111001"),
		("100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","101010011011","101010011011","101010011010","100010001010","100001010110","100101100101","100001010101","100101100110","011101000100","011101000101","100001010110","100001010110","100001010110","101010011010","100010001010","101010011010","101010011010","100001111001","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100010001010","100110001010","101010101100","101010011011","101010101100","100010001010","100101111000","100101100110","100001010101","011001010101","011001010101","011101000100","100001010110","100101100110","100101100110","101010011010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111000","100001111000"),
		("100001111001","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","100010001010","100001111000","100001111000","100001010110","100001010101","011101000101","011001010101","011001010101","100101100110","100001010110","100001010110","100101111000","100001111000","100010001010","100010001010","100110011011","100110011011","100110011011","100001111001","100001111000"),
		("100010001010","100001111001","100001111001","100001111000","100010001010","101010011011","101010011011","100110001001","100101111000","100101100111","011101000100","011101000100","011101000101","011001010101","011001010110","100001010110","100001010110","100010001010","100001111000","100001111000","100110001010","100110001001","100001111001","100110011011","100110011011","101010011010","100001111000"),
		("101010011011","100010001010","100001111001","100001111000","100001111000","101010011010","100110001010","100001111000","011000110100","100101100101","011100110011","011100110011","100001010110","010101000101","011001010110","100001010110","100101100111","100001111000","100001111000","100110001010","101010011010","100110001010","100001111001","100110001010","100110011011","100110001010","100001111001"),
		("101010011011","100110001010","100001111000","100001111000","100001100111","010100110011","010000100010","010000100010","010000100001","100001010110","011101000100","011101000100","011101000100","010101000101","011001010110","100001010110","100101111000","100001111000","100110001010","101010011010","101010011010","101010011010","100001111000","100001111000","100010001010","100001111000","100001111000"),
		("100110001001","011101010110","010100110100","010000100010","001100100001","001000100010","001000100001","001100100001","001100100001","100001100111","011101000100","011100110011","011101000100","011101100110","100001100111","100001010110","011101100110","100110001001","100110001010","100110001010","101010011010","101010011010","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("010000100010","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","100101111000","011101010110","011101000100","011101000100","100001111000","100101111000","100101111000","001100110011","001100110011","100110001001","100110001001","100110001010","100110001010","100110001010","100001111000","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010100110100","100001111000","100001111000","100001010110","100001000101","100101111000","100001100111","100110001001","001100110011","001100100010","001000100010","011101100110","100110001010","100110001010","100110001010","100001111000","100001111001","100110001001","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010101000101","100001111000","100110001001","100001010110","100001010110","011101010110","100001111000","100110001001","001100100010","001100100010","001000100010","001000100010","001100100010","100001111000","100001111000","100001111001","100110001001","100110001010","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001100110011","100001100111","100001111000","011001010110","100110001001","001100110011","001100100010","001000100010","001000100010","001100100010","001000100010","001100100010","100001111000","100001111000","100110001010","100110001010","100001111000"),
		("001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010110","010101000100","011001010110","011101100110","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010","001000100010","100001111000","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","011001010110","010101000100","010101000101","001000100010","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100010","100001111000","100001111001","100001111000","100001111000"),
		("001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100001111000","011001010110","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100001111000","100001111001","100110001001","100010001010"),
		("001000010001","001000010001","001000010001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","011001010110","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100101111000","100110001001","100001111001","100010001010"),
		("001100100001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","011101100110","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000010001","001000100010","001000100010","001000100010","100101111000","100110001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","010000110011","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100101111000","100010001010","100001111001","100001111001"),
		("001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","010000100010","010100110100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100110001001","100010001010","100010001010","100110001001"),
		("001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","010101000101","001100110011","010100110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100110001001","100110001001","100010001010","100110001001"),
		("001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","011001010110","001100110011","010100110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100110001001","100010001010","100110001001","100001111001"),
		("001000100001","000100010000","001000010001","001000010001","001000010001","000100010000","001000010001","001000010001","001000100010","001000100010","001000100010","010101000101","010101000101","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","100110001001","100110001001","100110001001","100110001001"),
		("001000100010","001000010001","001000010001","001000010001","000100010000","000100010000","001000010001","001000010001","001000100010","001000100010","001000100010","011001010110","010101000101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001100100010","100110001001","100110001001","100110001001","100110001001"),
		("001000100010","001000010001","100001100111","100001010101","011101000100","010000100010","011000110100","011000110011","001000100010","001000100010","001000100010","011001010110","011001010110","010100110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","010000110011","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","011101000101","100101100111","100001010101","011101000100","011100110011","001100010001","001000100001","001000100010","001000100010","001000100010","010101000100","011001010110","010100110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","011101100110","100110001001","100110001001","100110001001","100110001001"),
		("001100100010","100101100111","100001010110","011101000100","011000110100","001100010001","000100010000","000100010000","001000100010","001000100010","001000100010","001000100010","010101000101","010100110100","001000100010","001000010001","001000100010","001000100010","001000010001","001000010001","001000100010","001000100010","100001111000","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","100101100111","100001010101","011100110011","001000010001","000100010000","000100010000","000100010000","001000100001","001000100001","001000100010","010101000100","010101000100","010100110100","001000100010","001000010001","001000100010","001000100010","001000010001","001000010001","001000010001","001000010001","001000100010","100110001001","100110001001","100110001001","100110001001"),
		("010000110011","100101100110","011000110100","001100010001","001000010001","000100010000","000100010000","000100010000","000100010000","001000100010","001000100010","001100100010","001100100010","010100110100","001000100010","001000010001","001000100010","001000010001","001000010001","000100010000","001000010001","001000100001","001100100010","100101111000","100110001001","100110001001","100110001001"),
		("001000100010","010000100010","001000100010","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000100010","001000010001","001000100001","010100110100","001100100010","001000100001","001000100001","001000010001","000100010000","001000010001","001000010001","001000010001","001100100010","100001111000","100110001001","100110001001","100110001001"),
		("001000100001","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000100001","001000010001","001000100010","010000110011","001100100010","001000100001","001000010001","001000100001","000100010000","000100010000","000100010000","001000010001","001000010001","011001010110","100001111000","100001111000","100001111000"),
		("001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","011001010110","011001010110","010100110100","001100110011","001000100010","001000010001","001000100001","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","010100110100","100001100111","100001111000"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","010101000101","010101000101","010000110011","001100100010","001000100001","000100010000","001000010001","000100010000","000100010000","000100010000","000100010000","001000010001","010000100010","011000110011","011000110011","011000110011"))
	-- 0
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100110001001","100110001010","101010011011","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100010001010","100001111001","100010001001","101010011011","101010011011","101010101100","101010101100","101010011011","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","100110001010","100010001010","100110001010","100110011011","101010011100","101010101100","101010101100","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010101100","101010011011","100110001010","100010001010","100110011011","101010011011","101010001001","100101110111","101010001001","101010011011","101110101100","101010101100","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100110001010","100010001010","100110001001","100101110111","011101000011","011100110011","011101000011","011101000100","100001100110","101010011010","101010011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110011011","101010011011","100110001010","100110001010","100110001010","100110001010","100001100111","100101100101","100001010100","010100100010","010000100001","010000100001","010100100010","010100100010","011101000100","100101111001","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001011","100110001011","100110011011","100110001010","101010011011","101010101100","101010011011","100001010101","011100110011","011000110010","010100100001","010000100001","010000100001","010000100001","010000100001","010100100010","100001100111","101010011011","100110011011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","100110011011","101010011011","101110101100","101110101101","101010011011","100001010101","010100100010","011000110011","011000110011","011000110011","010100110011","010100100010","010100100010","010100100010","100001100111","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010101100","101110101101","101110101100","101110101100","101010011011","011101000100","011000110011","011101000101","100001010101","100101010110","100101100110","100101100110","100101100110","011101000100","100001100111","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011100","101110101101","101110101101","101110101100","101010001001","011000110011","011000110011","011101000101","100001000101","100001010110","100101100110","100101100110","100101100111","100001000101","100001111000","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010101100","101110101101","101110101101","101010101100","100101100111","011100110011","011101000100","011101000100","011100110100","011101000100","100001010110","100101010110","100101100110","100001010101","100110001001","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101101","101010011100","100110011011","100110011011","100110011011","101010101100","101110101101","101110101101","101010011011","100001000101","011101000100","011101000101","011101000101","011101000101","011101000100","100001010101","011101000100","011101000100","100101111000","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110001011","100110011011","101010011011","101010101100","101010101100","100001010110","011101000101","011101000101","011101000101","100001010101","011101000101","100001010110","100101100110","100001100110","100101111001","100110011010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100110011011","100110011011","100110001010","101010011011","101010101100","101010001010","100001010110","011101000100","011101000100","011101000101","011101000100","100001010101","100101100110","100101100111","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010","100110001001","100001100110","011101000100","011101000101","011101000100","100001000101","100001010110","100101010110","100101111000","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100001111000","100001100111","011101000101","011101000100","100001000101","011101000100","100001000101","100001010101","100101100111","100110001010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100010001010","100110001010","101010011011","100001111000","011101000100","100001010101","011101000100","011101000100","100001010101","100001100110","100001100110","100001100111","100110001010","101010011010","100110011010","101010011010","100110001010","100110001010","100110011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110011010","100010001001","100010001001","100001111001","100001100111","011001010101","010000100010","010000100010","011101000101","011100110100","011101000100","011101010101","011001010101","011101010110","100110001001","101010011011","101010011010","100110001010","100110001010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100010001010","100110001001","100001101000","011101010101","010100110011","001100100001","001100100001","001000100001","001100100010","011001010101","011101000100","011101000100","011101010101","011001010101","011101100110","100110001001","101010011010","100110001010","100001111000","100001111001","100010001001","100110001010","100110011010","101010011011","100110011010","100010001001","100001111000"),
		("011101100111","011001000100","010000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","011001010110","100001100111","100001000101","011001010101","010101000101","011101100110","100001110111","010101000101","100001101000","100001111001","100010001001","100110001010","100010001001","100001111001","100110011010","101010011011","100110001010","100001111001"),
		("001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","100001111000","100001010110","011001000100","010101000101","100001100111","100001111000","001100100010","001100100010","010101000101","100110001001","101010011011","100110001010","100001111001","100110001010","100110011011","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","011101100111","100110001010","100001111000","100001010110","011001010101","100001111000","011101101000","001100100010","001100100010","001000100010","010000110011","011101101000","100110001010","100001111001","100001111001","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100001","001100100010","001100100001","011001010101","100001111001","100001111001","100001100111","100001111000","100110001001","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","011101101000","100110001001","100001111000","100001111000","100001111000","100001111001"),
		("001000100010","001100100010","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001100100010","011001010101","011001010110","011101100111","100001111000","100001111000","010000110011","001100100010","001100100010","001100100010","001100100010","001000100010","011001010110","100110001010","100001111001","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010","010101000101","011101100111","011101100111","100001111000","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010110","100110001010","100001111001","100001111001","100010001001","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","010101000100","011101100111","011101100110","011001010110","010101000101","001100100010","001100100010","001100100010","001000100010","001100100010","001000100010","010101010101","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010001000100","011101100111","011001010110","011001010101","010101000101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010101","100110001001","100001111001","100110001001","100110001010","100001111001"),
		("001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010000110011","011101100110","011001010110","011001010101","010101000100","001100100010","001100100010","001000100010","001100100010","001100100010","001000100010","011001010101","100110001001","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010000110011","011101100110","011001010110","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001100100010","001000100010","011001010110","100110001001","100001111001","100001111001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","011101100110","011001010110","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100010001001","100001111000","100001111001","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","011001010110","011001010110","010101000101","010001000100","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","011101110111","100010001001","100110001001","100010001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001100110011","011001010110","011001010101","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001100110011","100001111000","100110001001","100110001001","100010001001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100001","001100110011","011001010110","011001010101","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100010001010","100010001001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100001","001100110011","011001010101","010101000101","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100110001001","100010001010","100010001001","100110001001"),
		("001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001100110011","011001010101","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001"),
		("001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001100100011","010101000100","010101000100","010101000100","010000110011","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100010001001","100110001001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","001000100010","001100100010","010101000100","010101000100","010000110100","001100110011","001000100010","001000100010","001000100010","001000100001","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100110001001","100001111000"),
		("001000010001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","000100010001","001000100001","001000100010","001100100010","010000110100","010000110100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","011101100110","100110001001","100110001001","100110001001","100010001001"),
		("000100010000","000100010001","000100010001","000100010000","000100010000","000100010001","000100010000","000100010000","001000100001","001000100010","001000100010","010000110011","010000110011","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001100100010","011001010110","100010001001","100110001001","100110001001"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000100010","001000100010","001100110011","010000110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000010001","001000010001","011001100110","100110001001","100110001001"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","000100010001","001000010001","001000100001","001000100010","010000110011","010000110011","001100110011","001000100001","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000100001","000100010000","000100010000","001000100010","011001010101","100110001001"),
		("000100010001","000100010001","000100010001","000100010001","001000010001","001000010001","000100010000","000100010000","000100010001","001000010001","010000110100","011001010110","010101010101","010000110011","001000100001","001100100010","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","001000100001","010101000101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010001","001000010001","010101000101","011101100111","011001010110","010101000100","010001000100","010000110011","001100100010","001000010001","001000010001","010001000100","001100110011","001000010001","000100010001","000100010000","001000010001","010000100010","010100110011"),
		("000100010001","000100010000","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010101000101","011101100111","011001010101","011001010101","011001010110","010000110011","001000100010","001000010001","001000010001","011001010110","100001111000","010101000101","001000100001","000100010000","001000010001","010000100010","011000110011"),
		("001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010101000101","011101100111","011001010101","011001010101","011001010110","010000110100","001100100010","001000100001","001000010001","011001010110","100010001001","100001111001","011101100111","010000110011","001000100001","001000010001","010000100010"),
		("001000010001","001000010001","000100010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010101000101","011001100110","010101010101","011001010101","011001010110","010001000100","001100100010","001000010001","001000010001","011101100110","100001111000","100001111000","100001111000","100001111000","011001010110","001100110010","001000100001"),
		("000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000100001","010101000100","010101010101","010101000100","010101000100","010101010101","010000110100","001000100001","000100010001","001000100001","011001010110","011101100111","011101100111","011101100111","011101100111","011101100111","011101100110","011001010110"))
	-- 1
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001100110","100001010101","100101100110","100001100110","100101111000","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100101111001","100001100101","011000110010","011000110010","010100110010","010100100010","011000110010","011101010101","100110001001","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001001","100101100110","100001000011","010100100010","010000100001","010000100001","010100100010","010100100010","010100100010","100001100110","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011100","101010011011","100001010101","011100110011","011000110010","010100100010","010000100001","010000100001","010000100001","010000100010","010100100010","011101010101","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100001010101","010100100010","010100110010","011000110011","011101000100","011101000100","011101000100","011101010101","011101000100","011101000101","101010011011","101010011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110011011","101010011011","100110001010","100110001010","100001010101","010100100010","011101000100","100001000101","100001010101","100101100111","100101100111","100101100111","100101010110","011101010101","100110001001","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001011","100110001011","100110011011","100110001010","101010011011","100001010110","011000100010","011101000100","011101000101","100001010101","100001010110","100101100111","100101100111","100101010110","100001010110","100101111001","100110001001","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","100110011011","101010011011","101010101100","100001100110","011000110011","011101000100","011101000100","011101000100","011101000100","100001010101","100001000101","100001010101","100101110111","100110001001","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010101100","101110101101","101010011011","100001010101","011100110011","011101000100","011101000100","011101000101","011101000100","100001010101","100001010101","100001010110","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101101","101010011100","100001010110","011101000100","011101000100","011101000101","100001010101","011101000100","100001010101","100101100110","100101100111","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101010101100","101010101100","100101111001","100001000101","011101000100","011101000100","011101000100","011101000100","100001010101","100101100110","100101100111","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101101","101010011100","100110011011","100110011011","100110011011","101010101100","101110101100","101010101100","101010011011","100001100110","011101000100","011101000101","011101000100","011101000100","100001010110","100101010110","100101111000","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110001010","100110001010","101010011011","101010101100","100110001010","100001010110","011101000100","011101000101","011101000100","011101000100","100001010101","100101100110","100001111000","100001111000","100010001001","100110011010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100110011011","100110001010","100110001010","100001111000","011001000100","011101000101","011101000100","011101000100","011101000100","011101000101","100001010110","100101111001","100110001010","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","100110011011","100110001010","011101100110","010000110010","001100100010","011001000101","011101000100","011101000100","011101000100","011101000101","100001100111","100110001010","101010011010","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100001111000","011101010110","010100110011","001100100010","001100100010","001100100010","010101000101","100001010110","100001000101","100001010101","100001010101","100101100111","100110001010","101010011010","101010011010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110001001","011101010110","010100110011","001100100010","001000100010","001100100010","001100100010","001100100010","001100110011","100001111000","100001010110","100001010101","011101010110","100001100111","100001110111","011101100111","100110001010","101010011010","101010011010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("011001000101","010000110011","001100100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100001111000","011101010101","011001000101","011101100111","011101100111","001100100010","010000110100","100001111000","100110001010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("001100100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100001","001000100010","001000100010","011001010110","100110001010","011101010110","011001000101","100001100111","011101100111","001100100010","001100100010","001100110011","011101111000","100010001010","100110001010","100110001010","101010011011","100110011010","100010001001","100001111000"),
		("001000100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","001100100010","010000110011","100001111000","011001010101","010101000100","100001100111","011001010110","001100100010","001100100010","001100100010","011001010110","100110001010","100010001001","100001111001","100110011010","101010011011","100110001010","100001111001"),
		("001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010","010101000101","011001010101","011001010101","011101100111","010000110100","001100100010","001100100010","001100100010","011001010110","101010011011","100110001010","100001111001","100110001010","100110011011","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","010101000100","011001010110","011001010110","011001010110","001100110011","001100100010","001100100010","001000100010","011101100110","101010001010","100110001010","100001111001","100001111001","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001000100010","001100100010","001100100010","001000100001","001000100001","001000100001","001000100001","001100100010","001000100010","010000110011","011101100110","100001111000","011101100110","010000110011","001100100010","001100100010","001100100010","100001111000","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111001"),
		("001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001100100010","001100100010","001100110011","011101100110","100001111000","011101100110","010000110011","001100100010","001100100010","010000110011","100110001001","100110001001","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001100100010","001100100010","011001010110","100001111000","011101100110","010000110011","001100100010","001000100010","010101000100","100110001001","100110001010","100110001010","100110001010","100001111001","100001111001","100010001001","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001100100010","001100100010","010101000100","011101100110","011001100110","010000110011","001100100010","001000100010","010101000101","100110001010","100110001010","100110001001","100001111001","100001111001","100010001001","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","010000110100","011001010101","011001010110","010000110011","001100100010","001000100010","010000110100","100110001001","100110001010","100001111001","100001111001","100001111001","100110001001","100110001010","100001111001"),
		("001000100001","001000100001","001000100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","010000110011","011001010101","011001010110","010000110011","001000100010","001000100010","010000110100","100110001001","100001111001","100001111000","100010001001","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001100110011","011001010101","011001010101","010000110011","001000100010","001000100010","010000110100","100001111001","100001111001","100110001001","100110001001","100001111001","100001111001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","000100010001","001000010001","000100010001","000100010001","001000010001","001000100010","001100100010","010101000101","011001010101","010000110011","001000100010","001000100010","010001000100","100001111001","100110001001","100110001001","100001111001","100001111000","100001111001","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","000100010001","000100010001","000100010000","000100010000","001000010001","001000100010","001100100010","010101000101","010101000100","001100100010","001000100001","001000100010","010101000100","100001111001","100001111001","100001111001","100010001001","100110001001","100010001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010001","001000100001","001100100010","010101000101","010000110100","001000100001","001000100001","001000100010","010101000101","100001111001","100001111000","100001111000","100110001001","100110001001","100010001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001000010001","001100100010","010101000100","010000110011","001000100001","001000100001","001000100010","010000110011","100001111000","100001111001","100110001001","100110001001","100110001001","100010001010","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001100100010","010101000100","010000110011","001000100001","001000100001","001000100010","001000100010","010001000100","100001111000","100110001001","100110001001","100110001001","100010001010","100010001001","100110001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010001","001100100010","010000110100","010000110011","001000100010","001000100001","001000100010","001000100010","001000010001","010000110011","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001100100010","010000110100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000101","100001111000","100110001001","100110001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001100100010","010000110011","001000100001","001000100001","001000100010","001000100010","001000100001","001000100010","001000100010","001000010001","001100110011","100001111000","100110001001","100010001001","100010001001"),
		("001000100001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000100010","010000110100","001100100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000010001","001000010001","010101000100","100101111000","100101111001","100101111001"),
		("001000010001","000100010000","000100010001","000100010000","000100010000","000100010001","000100010000","000100010001","001000010001","000100010000","000100010000","000100010000","001000100001","010101000100","010000110100","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000010001","001100100010","011001000100","100001010101","100001010110","100001100110"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","001000100001","010101000100","011001010101","010000110100","001000100010","001000100010","001000100001","001100100010","001100110011","001000010001","001100100010","010100100011","011000110011","011000110011","011101000100"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","000100010001","001000010001","000100010000","000100010000","000100010000","001000100001","010101000100","011001010110","011001010110","001100110011","001000100010","001000010001","001100110011","100001111000","010101000101","001100100010","011000110100","011001000100","011000110011","011000110011"),
		("000100010001","000100010001","000100010001","000100010001","001000010001","001000010001","000100010000","000100010000","001000010001","000100010001","000100010000","000100010000","001000100001","010101000100","011001010110","011001010110","010001000100","001000100010","001000010001","001100100010","100001111000","100110001001","100001111000","100001111000","100101111001","100001100111","011101010101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001000100001","010000110100","011001010110","011101100110","010101000101","001000100001","000100010001","001100110011","100001111001","100110001001","100110001001","100110001001","100110001001","100110001001","100101111001"),
		("000100010001","000100010000","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001000100001","010000110100","011001010110","011101100110","010101010101","001000100001","000100010001","010001000100","100010001001","100010001001","100110001001","100110001001","100110001001","100110001001","100110001001"),
		("001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","000100010000","000100010000","001000100010","010101000100","011001010110","011101100110","010101000101","001000100001","000100010000","010101000101","100001111001","100001111001","100001111001","100001111001","100010001001","100010001001","100001111001"),
		("001000010001","001000010001","000100010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","000100010000","000100010000","001000100001","010101010101","011001010110","011001010110","010101000101","001000100001","000100010000","010101000101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000100001","010101000100","010101010101","011001010101","010101010101","001000100010","000100010001","010101000100","011101100111","011101100111","011101100111","011101100111","011101100111","011101100111","011101100111"))
	-- 2
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100001111001","100101111001","100101111000","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011010","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011100","100110001001","100101100110","100101100101","100001000100","011101000100","011101000100","100101100111","101010011011","101010101100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","100110001010","100101010101","011101000011","011000110010","010100100010","010100100010","010100100010","011000110011","100001100111","101010011011","101010011100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100101100111","011000110010","010000100001","010100100010","010100100010","010100100010","010000100010","010100100010","011001000100","101010011011","101010101100","101010011100","101010011011","100110011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110011011","100110001001","100101010101","011000110010","010000100001","010000100001","010000100001","010100110011","011101000100","011101010101","011000110011","100110001001","101010101100","101010011011","100110001001","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001011","100110011011","100101111000","011101000011","010100100010","011000110011","011101000100","100001010101","100001010110","100101100111","100101100111","011101000101","100001100111","101010011011","100110011010","100110001001","100110001001","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","100110001001","011000110011","011000110011","100001010101","100001010101","100101100110","100101100110","100101100111","100101010111","100001010110","100001111000","100110001010","100110001001","100110001001","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011011","011101000101","011000110011","011101000101","011101000101","100001010101","100001010110","100001010110","100001010101","100001010110","100101111000","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","100101111000","011000110011","011101000100","011101000100","011101000100","011101000101","100001010101","100001010101","100001010110","100101100111","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101010001010","011101000100","011101000100","011101000101","011101000100","011101000100","100101010110","100101100111","100101010110","100101100111","100110001010","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101101","101010011100","100110011011","100110011011","100110011011","101010101100","100110001001","011101000100","011101000100","011101000101","011101000101","011101000100","100001010101","100101100110","100101010110","100101111000","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110001010","100110001010","100110001010","100001010110","011101000100","011101000100","011101000101","011101000100","100001010110","100101010110","100101010110","100101111001","100001111001","100001111000","100010001001","100110011010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100110011010","100110001010","100110001010","100110001010","100001100111","011101000100","011101000100","011101000100","100001000101","100001010110","100101100110","100110001010","100110001010","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","100110011011","100110011010","100010001001","100110001001","100001100111","011101000100","011101000100","011101000100","100001010101","100101010110","100101100111","100110001010","101010011010","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100010001001","100001111001","100110001010","100110001001","100010001001","100001100111","011101000101","011101000100","011101000100","011101000100","011101000101","100001010101","100101100111","100110001010","101010011010","101010011010","100110011010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110001010","100001111001","100010001001","100010001001","100010001001","100110001001","010101000100","010000110011","011101000101","011101000100","011101000100","100001010110","100001100111","100001100111","100001111000","010101000101","011101100111","100110001010","101010011011","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100001111001","100001100111","010101000100","001100100010","001100100010","011101010110","100001010110","011101000101","011001010101","011001010101","011101010110","100001111000","010000110011","001100100010","010001000100","100001111000","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100001111001","100001111001","100101111000","011101010110","010000100010","001100100001","001100100001","001000100010","010000110100","100001111000","100001010110","011001010101","011001010101","011001010110","100001111001","010101000100","001100100010","001100100010","010000110100","100001111001","100110001010","100110001010","101010011011","100110011010","100010001001","100001111000"),
		("100001111001","100001111001","100001100111","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","011101100111","100001111000","011001000101","011001010101","011001010110","100110001001","010101000100","001100100010","001100100010","001100110011","100001111001","100010001001","100001111001","100110011010","101010011011","100110001010","100001111001"),
		("100101111001","011101010101","010000100011","001000100010","001000100010","001000100010","001100100010","001100100010","001000100010","001000100010","011001010110","100001111000","011001000101","011001010101","100001111000","100110001001","010000110100","001100100010","001100100010","010000110011","100110001010","100110001010","100001111001","100110001010","100110011011","100110001010","100001111001"),
		("010000110011","001100100010","001000100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001000100010","010000110011","100001111000","011101100110","011001010110","011101100111","011101100111","001100110011","001100100010","001000100010","010101000100","100110001010","100110001010","100001111001","100001111001","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","010101000101","011101100111","011101100111","011001010110","011001010110","001100110011","001100100010","001100100010","010101000101","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111001"),
		("001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","010000110011","100001100111","011101100111","011001010110","011001010110","010000110011","001100100010","001100100010","010101000101","100110001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100001100111","011001010110","011001010110","010000110100","001100100010","001000100010","010101010101","100110001010","100110001010","100110001010","100001111001","100001111001","100010001001","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001100100010","001100100010","001100100010","001100100010","010101000100","011101100110","011001010110","011001010110","010001000100","001100100010","001000100010","011001010110","100110001010","100110001001","100001111001","100001111001","100010001001","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","001000100010","001100100010","001100100010","001100100010","001000100010","010000110011","011001010110","011001010110","011001010110","010101000100","001000100010","001000100010","010101010101","100110001010","100001111001","100001111001","100001111001","100110001001","100110001010","100001111001"),
		("001000100001","001000100001","001000100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000100010","001100100010","001000100010","001000100010","010000110011","011001010110","011001010110","011001010110","010101000100","001000100010","001000100010","011001010110","100010001001","100001111000","100010001001","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100010","001100100010","001000100010","001000100010","010000110011","010101010101","011001010110","011001010110","010001000100","001000100010","001000100010","011001010110","100001111001","100110001001","100110001001","100001111001","100001111001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","010000110011","010000110011","011001010101","011001010101","010000110011","001000100010","001000100010","011101100111","100110001001","100110001001","100001111001","100001111000","100001111001","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","000100010001","000100010001","000100010000","001000100001","001000100010","001000100010","010000110011","001100110011","010101010101","011001010101","010000110011","001000100010","001100100010","011101100111","100110001001","100001111001","100010001001","100110001001","100010001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010001","001000100010","001000100010","010000110011","001100100011","010101000100","010101010101","001100110011","001000100010","001100100010","011101101000","100001111000","100001111000","100110001001","100110001001","100010001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000010001","001000100010","001100110011","001100100011","010000110011","010101000101","001100100010","001000100010","001100100010","100001111000","100001111001","100110001001","100110001001","100110001001","100010001010","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","001000010001","001100110011","001100110011","001100100011","010101000100","001100100010","001000100001","001000100010","011101010110","100110001001","100110001001","100110001001","100110001001","100010001010","100010001001","100110001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000010001","001100110011","001100100011","001100100010","010000110011","001000100010","001000100010","001000100001","001100100010","100101111000","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001100110010","001100100011","001000100010","001100100010","001000100001","001000100001","001000100010","001000100010","011001010101","100110001001","100110001001","100010001001","100110001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001100100010","001100100010","001000100001","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001100100010","001100100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","011001010110","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","000100010000","000100010001","000100010000","000100010000","000100010001","000100010000","000100010001","001000010001","001000010001","001000010001","000100010000","001100100010","001000100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100001","001000010001","010000110011","011101000101","100001100110","100001100111","100101111000","100110001001"),
		("001000100001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000100001","001000010001","000100010000","001100100010","001000100001","001000010001","001000100001","001000100001","001000100010","001000100001","001000100001","001000100001","010000100010","011000110011","011000110100","100001010101","100001010101","100001110111"),
		("001000100010","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","000100010001","001000010001","000100010000","000100010000","000100010001","001100100010","001000100001","000100010000","001000100001","001000100001","001000100001","001000100001","001000100001","000100010001","010000100010","010100100010","010100100010","011000110011","011101000100","011101000101"),
		("001100100010","000100010001","000100010001","000100010001","001000010001","001000010001","000100010000","000100010000","001000010001","000100010001","000100010000","000100010000","001100110010","001000100001","000100010000","001000010001","001000100010","001000100001","001000100010","011001010110","010000110011","011001010110","100001100111","011000110100","010100100010","011000110011","011101000100"),
		("001100100010","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","001000010001","000100010000","000100010000","001100100010","001000100001","000100010000","000100010000","001000100010","001000100001","001000100010","100001111000","100010001001","100110001001","100110001001","100001111000","011001000100","011101000100","100001100111"),
		("001100100010","000100010000","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001100100010","001000100001","000100010000","000100010000","001000100001","001000100001","001100110010","100001111000","100010001001","100010001001","100110001001","100110001001","100001111000","100001111001","100110001001"),
		("001000100010","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","000100010000","000100010000","000100010001","000100010000","000100010000","001100100010","001000100001","000100010000","000100010000","001000010001","001000010001","010001000100","100001111001","100001111000","100001111001","100001111001","100001111001","100010001001","100010001001","100001111001"),
		("001000100001","001000010001","000100010001","000100010001","000100010000","000100010001","001000010001","000100010001","000100010000","000100010000","001000010001","000100010001","001100100010","001000100001","000100010000","000100010000","001000010001","001000010001","010101000101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","001000100010","001000100001","000100010001","000100010000","001000100010","001000100010","010101000100","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111","011101100111","011101100111"))
	-- 3
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011010","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001001","100110001001","100110001001","100101111001","100001111001","100110001010","101010011011","101010011011","101010011100","101010101100","101010011100","101010011100","101010011011","100110011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001011","100101111001","100101110111","100101010101","100001010100","011101000100","100001010100","100001010101","100001100111","100110001001","101010011011","101010101100","101010101100","101010011100","101010011011","100110001001","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001001","100101010101","011101000011","011000110010","010100100010","010100100010","011000110011","011000110011","011000110100","100001111000","100110011010","101010011011","101010101100","101010011011","100110011010","100010001001","100110001001","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100001100110","011000110011","011000110010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","100001100110","100110001001","100110001010","101010011011","100110001010","100110001001","100110001001","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100001010110","010100100010","010000100001","010000100001","010100100010","011000110011","100001010101","100001010101","010100100010","011001000100","100110001001","100010001010","100110001001","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100101100111","011000110011","010100110010","011000110011","011101000101","100101010110","100101100111","100101100111","011101000100","011000110100","100110001010","100110001010","100110001010","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100101110111","011101000100","100001010101","100001010101","100001010110","100001010110","100101100111","100101100111","100001010110","011001000100","100110001001","100110001001","100110001001","100110001010","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100101111001","011101000100","011101000101","011101010101","100001010101","100001010101","100001010101","100001010110","100001010110","011101000101","100101100111","100001111001","100110001001","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110001010","100001010110","011101000100","011000110011","011101000100","100001010101","011101000101","100001010101","100101010110","100001010110","100101100111","100110001001","100110001001","100001111001","100001111000","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100101111001","100001010101","011000110100","011101000100","100001010110","100101010110","100101010111","100101010111","100101010110","100101100111","101010011010","101010011010","100110001010","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","100110001001","100001100110","011101000100","011101000100","100001010101","100001010111","100001010111","100101010111","100101100111","100110001001","100110011010","100110001010","101010011010","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001001","100110001010","100101100111","011101000101","011101000100","011101000101","100001010110","100001010110","100101010110","100101100111","101010011010","101010011011","101010011010","101010011010","100110011010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110001010","100010001001","100010001001","100010001001","100010001001","100001010110","011101000100","011101000100","100001010101","100001010110","100001010110","100001010110","100001111000","100110001010","101010011010","101010011010","101010011010","101010011010","101010011011","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100001111001","100110001010","100110001010","011101000101","011101000100","100001000101","100001010110","100001010110","011001010101","011001010101","011101100111","100001111000","011101100111","100001111000","100001111000","100110001001","100010001001","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100001111001","100001111000","100001111000","100110001001","101010011011","100110001001","011101010101","011101000100","011101000100","100001000101","100001010101","011001010101","011001010101","011101010110","001100100011","001100100010","001100100010","001100100010","010000110011","010000110100","011101101000","100110011010","101010011011","100110011010","100010001001","100001111000"),
		("100001111001","100001111000","100001111000","100001111000","100110001010","101010011010","011001000101","011001000100","011000110011","011000110011","011000110011","011101000101","011001010101","011001010101","100001111000","010000110100","001100100010","001100100010","001100100010","001100100010","001100100010","010000110100","100001111001","100110011010","101010011011","100110001010","100001111001"),
		("101010011011","100110001001","100001111000","100001111001","100110001001","011101010110","001100100010","011001000101","011101000100","011000110011","011100110100","011101000101","011001000101","011001010101","100001111000","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101101000","100110001010","100110011011","100110001010","100001111001"),
		("101010011011","100110001001","100001111001","100001111000","011001000101","001100100010","001000100010","010000110100","100001110111","011101010101","011101000100","100001000101","011001010101","011001010110","100110001001","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010110","100001111001","100010001001","100001111001","100001111000"),
		("101010011010","100110001001","100001100111","010100110100","001100100010","001100100010","001100100010","001100100010","011101100110","100001111000","100001100110","100001010110","011101010110","100001111000","100110001010","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010101","100001111001","100001111000","100001111000","100001111001"),
		("101010001010","100001100110","010000110011","001000100001","001000100001","001000100010","001000100010","001100100010","010101000101","100001111001","100010001010","100001111001","100001100111","100001111000","100110001001","010101010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010101","100001111001","100001111000","100001111000","100001111000"),
		("011001010101","001100100010","001000100001","001000100010","001000100010","001000100001","001000100010","001000100010","001100110011","011101100111","100001111001","011101100111","100001111000","100001100111","011101100111","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010101000101","100001111001","100001111001","100010001001","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010101","011001010110","011001010110","011101100110","011001010110","011001010101","001100110011","001100100010","001100100010","001100100010","001100100010","001100100010","010101000101","100001111001","100010001001","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001000100010","010101000100","011001010110","011001010101","011001010101","011101100110","011001010110","001100110011","001000100010","001100100010","001100100010","001100100010","001100100010","011001010101","100010001001","100110001001","100110001010","100001111001"),
		("001000100001","001000100001","001000100010","001000100001","001000100010","001100100010","001100100010","001000100010","001000100010","001100100010","001100110011","011001010110","011001010101","011001010101","011001010110","011001010110","010000110011","001000100010","001100100010","001100100010","001100100010","001100100010","011101100111","100010001001","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","011001010101","011001010101","011001010110","011001010110","010000110100","001000100010","001100100010","001100100010","001100100010","001100100010","011101100111","100010001001","100001111001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010101","011001010110","011001010110","011001010110","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100110011","100001111000","100010001001","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","010101000101","011001010110","011001010110","011001010110","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","100001111000","100010001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010101","011001010110","011001010101","010000110100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","011101100111","100110001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000100010","001100100010","001000100010","001000100010","001000100010","001100110011","011001010101","011001010110","011001010101","010000110100","001100100010","001000100010","001100100010","001000100010","001000100010","001000100010","011001010110","100110001010","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100001","001100110011","011001010101","011001010110","010101010101","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","010101000101","100110001010","100010001001","100110001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000100001","001000100010","001000100010","001000100001","001100110011","010101000101","011001010101","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","011101100111","100110001010","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010001","001000100001","001000100010","001000100010","001100110011","010000110011","011001010101","010101000100","010000110100","001100110011","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","010000110011","100001111000","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010000","001000010001","001000100010","001000100010","001100110011","001100110011","010101000100","010101000100","010000110011","001100100010","001000100001","001000100010","001000100010","001000100001","001000010001","001000010001","001000100010","100001111000","100110001001"),
		("001000100001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","001000010001","001000100010","001100110011","001100100010","010001000100","010101000100","010000110100","001100100010","001000100001","001000100001","001000100010","001000100001","000100010001","001000100001","001100100010","011101100111","100110001001"),
		("001000010001","000100010000","000100010001","000100010000","000100010000","000100010001","000100010000","000100010001","001000010001","000100010000","001000010001","001000100001","001100110011","001100100010","010000110011","010101000100","010000110100","001100100010","001000100001","001000100001","001000100010","001000010001","000100010000","001100100010","011001000100","011101000101","100001010110"),
		("001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001100110011","001100100011","001100100010","010000110100","010000110011","001100100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100001","011000110100","011000110100","011000110011"),
		("001000010001","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","000100010001","001000010001","000100010000","000100010000","000100010001","001100100010","001100100010","001000100010","010000110011","010000110011","001100100010","001000010001","001000100001","001000100001","001100110010","011101100110","001100100010","010000100010","011101000100","011101000100"),
		("001000010001","000100010001","000100010001","000100010001","001000010001","001000010001","000100010000","000100010000","001000010001","000100010001","000100010000","000100010000","001100100010","001100100010","001000100010","001000100001","001100100010","001100100010","001000010001","001000100001","001000100001","001100100010","100001111000","100001100111","010000100010","011000110011","100001010110"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","001000010001","000100010000","000100010000","001100100010","001100100010","001000100001","001000100010","010001000100","010000110100","001000100001","001000010001","001000100001","001100100010","100001111000","100110001001","011101010110","011001000100","011101010110"),
		("001000010001","000100010000","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001100100010","001000100001","001000010001","001100110011","011001010101","010101010101","010000110011","001000100010","001000100001","001000100010","011101110111","100110001001","100110001001","100001111000","100001111000"),
		("001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","000100010001","000100010000","000100010001","000100010000","000100010000","001100100010","001000100001","000100010000","001100100010","011001010101","011001010110","010101000101","001100110011","001000010001","001000100010","011101100111","100010001001","100010001001","100010001001","100010001001"),
		("001000010001","001000010001","000100010001","000100010001","000100010000","000100010001","001000010001","000100010001","000100010000","000100010001","000100010001","000100010000","001100100010","001000100001","000100010000","001000010001","010101000101","011001010110","010101000101","010000110011","001000100001","001000100001","011001010110","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000100010","001000100001","000100010001","000100010000","010000110011","010101010101","010101000100","010000110011","001000100010","001000100001","010101000101","011101100111","011101100111","011101100111","011101100111"))
	-- 4
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001001","100001111001","100001111001","100110001010","101010011011","101010011011","101010011100","101010101100","101010011100","101010011100","101010011011","100110011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001010","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011100","101010011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100101111000","100101100111","100101100110","100001100110","100101110111","100101110111","100101111000","100110001001","100110001010","101010011011","101010101100","101010011011","100110011010","100010001001","100110001001","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100101110111","100001010100","011100110011","011000110010","011000100010","011100110011","011101000011","011101000100","100001111000","100110001001","100110001010","101010011011","100110001010","100110001001","100110001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100101111000","100001000100","011100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011001000101","100110001001","100010001010","100110001001","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100101110111","011000110011","010000100001","010000100010","010100100010","010100110011","011001000100","011000110100","010100100010","011000110011","100110001010","100110001010","100110001010","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100101111000","011101000011","010100110010","011000110011","011101000101","100001010110","100101100111","100101100110","011000110011","010100100010","100101111000","100110001010","100110001001","100110001010","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110001001","100001010101","011101000101","100001010101","100001010101","100001010110","100101100111","100101100111","011101000101","010100110011","100001100111","100010001001","100110001001","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110001010","100001010110","100001010101","100001010101","100001010101","100001010101","100001010110","100001010110","100001010110","011000110011","100001100111","100110001001","100110001001","100001111001","100001111000","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100101100111","011101000101","011000110100","011101000100","100001010101","011101000100","100001010110","100101010111","011101000101","100001010110","100110001010","101010011010","100110001010","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","100110001001","011101010101","011000110011","011101000100","100101010110","100001010110","100001010111","100101010111","100101010110","100001010110","100110001010","100110011010","101010011010","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001001","100110001010","100001010110","011101000100","011101000100","100001010110","100001010110","100001010110","100101010111","100001010110","100101111000","101010011011","101010011010","101010011010","100110011010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110011010","100010001001","100010001001","100010001001","100001100110","011101000100","011101000100","100001010101","100001010110","100001010110","100001010110","100001010110","100101111000","100110001010","100110011010","100110001010","100110011010","100110011010","101010011010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100001111001","100101111001","011101000101","011101000100","011101000101","100001010110","100001010110","100001010110","011001010101","011001010101","100101111001","101010011010","101010011010","100110001010","100110001010","100110001010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100001111001","100001111000","100001111000","100110001010","101010011011","100001100111","011101000100","011101000100","100001010101","100001010110","100001010110","011001010101","011001010101","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001","100110001001","100110001010","101010011011","100110011010","100010001001","100001111000"),
		("100001111001","100001111000","100001111000","100001111000","100110001001","101010011011","101010011010","100001010101","011101000100","100001000101","100001010101","100001010110","011001000101","011001010101","011001010110","011001010101","011001010110","011001010110","011001010110","011001010110","011001010110","011101100110","011101101000","100110001010","101010011011","100110001010","100001111001"),
		("101010011011","100110001001","100001111000","100001111000","100001111001","100110001010","100110001010","100001010110","011000110011","011000110011","011101000100","100001010101","011001000101","011001010101","011101100111","001100100011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100011","011001010110","100110011010","100110001010","100001111001"),
		("101010011011","100110001001","100001111000","100001111000","100001111001","100001111001","100001100111","011101000101","011000110011","011000110011","011101000100","100001010101","011001010101","011001010110","100001111001","010001000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100001111001","100001111000"),
		("101010011010","100110001001","100001111000","100001111000","100001111001","011101100111","010000110011","011001000101","011101000101","011000110011","011101000100","100001000101","011101010110","100001110111","100110001001","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010101000100","100001111001","100001111001"),
		("101010011010","100110001001","100001111000","100001111000","011001010101","001100100010","001000100010","010001000100","100001111000","011101000101","011101000100","100001010101","100001100111","100001111000","100110001001","010101010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","010000110011","100001111001","100001111000"),
		("101010011010","100110001001","100001100111","010100110100","001100100010","001000100001","001000100001","001100100010","011101100111","100001111001","100001010111","100001010110","100001100111","100001111000","100110001001","010101000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100001111001"),
		("101010001010","011101010110","010000100010","001000100001","001000100010","001000100010","001000100010","001000100010","011001010110","100001111001","100001111001","011101100111","011101100110","011101100111","100001111000","010001000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","010000110100","100001111001"),
		("011001000101","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110100","011101100110","010101010101","010101000101","010101000101","011001010101","011001010110","010001000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","100001111000"),
		("001000100001","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","010101000100","011001010101","011001010101","011001010101","011001010110","010101000100","001100100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","010000110011"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","011001010101","011001010101","011001010101","011001010110","010101000100","001100100010","001000100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001"),
		("001000100001","001000100001","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010101","010101010101","010101010101","011001010101","010101000100","001100110011","001000100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001100100010","010101000101","010101010101","011001010101","010101010101","010101000100","010000110011","001000100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000010001","001000100001","001000100001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","010001000100","010101000101","011001010101","010101010101","010101000100","010000110011","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000010001","001000100001","001000100001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100001","001000100010","001100110011","010101000101","011001010101","010101000101","010001000100","010000110011","001100100010","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000010001","001000010001","001000100001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001100100010","010101000100","011001010101","010101000100","010001000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000100010","001000100010","001000100010","010000110100","010101000101","010001000100","010000110100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000010001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001000100010","001100110011","010101000101","010001000100","010000110100","010000110100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","010000110100","001000100010"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001100110011","010101000100","010001000100","010000110100","010000110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001"),
		("001000100001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001100110011","010101000100","010000110100","010000110100","010000110011","010000110011","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000010001","001000100001","010000110011"),
		("001000010001","000100010001","000100010001","000100010000","000100010000","000100010001","000100010000","000100010001","001000010001","001000010001","001000100001","001000100001","001100110011","010000110011","010000110100","010000110011","010000110011","010000110011","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","011000110100","011000110011"),
		("001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","001000010001","000100010001","001000010001","001000100001","001100110011","001100110011","010000110011","010000110100","010000110011","010000110011","001100100010","001000100001","001000100010","001000100010","001000100001","001100100010","001100100010","011000110011","011000110011"),
		("001000010001","000100010000","000100010000","000100010000","000100010000","001000010001","001000100001","000100010001","001000010001","000100010000","001000010001","001000010001","001100110010","001100100011","010000110011","010001000100","010000110100","010000110011","001100100010","001000100001","001000100001","001000100010","001000100001","001000010001","001000010001","010100110011","011101000101"),
		("001000010001","000100010001","000100010001","000100010001","001100100010","001000100001","001000100010","001000100001","001000010001","000100010001","000100010000","001000010001","001100110011","001100100010","001100100011","010000110011","010000110011","010000110011","001100100010","001000100001","001000100001","001000100010","001000100001","000100010000","001000100001","011000110100","011101000101"),
		("001000010001","001000010001","001000010001","001000010001","011001000101","001100110010","000100010000","001000100001","001000010001","001000010001","000100010000","001000010001","001100110011","001100100010","001100100010","001100110011","001100100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","000100010000","001000010001","001100100010","010100110011"),
		("001000010001","000100010001","001000010001","000100010001","001000100010","001100100010","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001100100010","001100100010","001000100010","001000100010","001100100010","001100100010","010000110011","010000110011","001100100010","001000100010","001000100001","000100010001","000100010001","001000100001","001000100010"),
		("001100100010","001000100001","001000010001","000100010000","001000010001","001000100001","000100010000","000100010000","001000010001","001000010001","000100010000","000100010000","001100100010","001100100010","001000100010","010001000100","010101000101","010101010101","011001010101","010101000101","010000110011","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010"),
		("001100100010","001000010001","000100010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","000100010000","000100010000","001100100010","001000100010","001000100010","010101010101","011001010110","011001010101","011001010101","010101010101","010000110100","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("001000100001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000100010","001000100001","001000010001","010001000100","011001010101","010101000101","010101000101","010101000101","010000110100","001100100011","001000100001","001000100010","001000100010","001000100010","001000100010"))
	-- 5
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011100","101010101100","101010011100","101010011100","101010011100","101010011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001001","100110001010","100110001001","100001111001","100110001001","101010011011","101010101100","101010101100","101010101100","101010011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","101010011010","100110001001","100110001001","100110011010","101010011011","101010101100","101010011011","100110011010","100110001001","100110001010","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011100","101010001001","100101110111","100001010101","100001010101","100001010110","100101110111","100110001010","101010011011","100110001010","100110001001","100110001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101010101100","100101111000","100001010100","011101000011","010100100010","010100100010","011000110010","011101000011","011101010101","100101111001","100110001001","100110011010","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101010011011","100001010100","011000110010","010100100010","010100100010","010000100010","010100100010","010100100010","010100100010","011101010110","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101010001010","011101000100","010100100010","010100100010","010100110010","011000110100","011101000100","011101000100","010100100010","011001000100","101010011010","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101010001001","100001010100","011101000100","011101000100","100001010101","100101100110","100101100111","100101100111","011000110100","010100110011","100101111001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110011011","100101111000","100001000101","100001010101","100001010101","100001010110","100101010110","100101100111","100101100111","100001000101","011000110011","100001111000","100001111001","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110011011","100101111000","011101000101","100001000101","011101000100","100001010101","100001010110","100001010101","100001010110","100001010110","011001000100","100110001001","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010101100","100110001010","100110001010","101010011011","101010011011","100110001010","100001100110","011101000100","011000110100","011101000100","100001010110","011101000101","100001010110","100101010110","011101000101","100110001001","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100101111000","100001010101","011101000100","011101000101","100101010111","100001010110","100101010111","100101010111","100001010110","100101111000","101010011010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110011010","100010001001","100110001001","100110001001","100110001010","101010011011","100101111000","100001010101","011101000100","011101000100","100001010110","100001010110","100101100111","100001100111","100001010111","100110001001","101010011010","100110011010","101010011010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100110001010","100110011010","101010101100","100110001001","100001010110","011101000100","011101000100","100001010101","100001010110","011001010101","011101010110","100101111000","101010011010","100110011010","100110001010","100110001010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100010001001","100010001001","100001111001","100001111001","100110001010","101010011011","101010101100","101010011010","100001100111","011101000100","011100110011","011101000100","011101010101","011001010101","011101010110","100110001001","101010011010","100110001010","100001111000","100001111000","100001111000","100010001001","100110001010","101010011011","100110011010","100010001001","100001111000"),
		("100010001001","100001111000","100001111001","100001111000","100110001010","101010011011","101010011011","100110001010","100001111000","100001010110","011101000100","011101000101","011101010101","010101000101","011101010110","100101111001","100110001010","100110001001","100001111000","100001111001","100110001001","100001111000","100001111001","100110001010","101010011011","100110001010","100001111001"),
		("101010011011","100110001001","100001111001","100001111001","100001111001","100110011010","100110001010","100001111000","100001111001","100001110111","011101000100","011101000100","011001010101","010101000101","011101010110","100101100111","100001111000","100001111000","100001111001","100110001010","101010011010","100110001001","100001111000","100010001001","100110011010","100110001010","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100010001001","100001111001","100001111001","100001111000","100110001001","100101111000","011100110100","011100110011","011101010101","011001010101","011101010110","100001010111","011101010110","010000110011","011001010101","011101100111","100001111000","100110001001","100001111000","100001111001","100110001010","100001111001","100001111000"),
		("101010011011","100110001010","100001111001","100001111000","100001111001","100001111000","100001111000","100110001001","100110001010","100101111000","011101000100","011100110100","011101000101","011101100111","100001100110","100001010110","100001111000","001100110011","001100100010","001100100010","001100100010","010000110011","010101000100","010101000101","011101100110","100001111000","100001111001"),
		("101010011011","100110001010","100001111000","100001111001","100110001001","100110001010","100001111001","100110001001","100001111000","100001100111","011101000100","011101000100","011101000101","100001111000","011101010110","100001100111","100010001001","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001100100010","001100110011","011001010110"),
		("101010011010","100110001001","100001111001","100010001001","100110001010","101010011010","100101111000","011001000101","010100110011","100001100111","100001100111","011101000100","100001010110","100001111000","011101010110","100001111001","100001111001","001100110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100110011"),
		("101010011011","100110001001","100010001001","100110001001","100110001001","100001100111","010100110011","001100100010","001100100010","011101100111","100010001001","100001100111","011101010101","011101100111","100001111000","100110001010","011101100111","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","100110001010","100110001001","100001111000","011101000101","010000100010","001000100010","001000100010","001000100010","011101010110","100001111000","100001111001","011101100110","011001010101","100001111000","100110001010","011001010101","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010"),
		("101010011011","100110001001","011101010110","010100110011","001100100010","001000100010","001000100010","001000100010","001000100010","010000110100","010101000101","010101000101","010101000101","010101010101","011001010101","011101100111","010101000100","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100101111000","010000110011","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","010101010101","010101010101","010101010101","011001010101","010001000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100001111000","001100100010","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101010101","010101010101","011001010101","011001010101","010101000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001"),
		("100110001001","100001111000","001100100010","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","010101010101","010101000101","010101000101","010101000101","010101000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001001","011101100111","001100100010","001000010001","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001100110011","010101000101","010101000101","010101000101","010101000100","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001010","011101100111","001000100010","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100001","001000100010","001100100010","010101000100","010101000101","010101000100","010101000100","010001000100","001100100010","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001"),
		("100110001010","011001010110","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","010000110100","010101000101","010101000100","010000110100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001"),
		("100110001001","011001010110","001000100001","001000010001","001000010001","001000010001","001000010001","000100010000","001000100001","001000100010","001000100010","001000100001","010000110011","010101000101","010101000100","010001000100","010001000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000010001"),
		("100110001001","011001010110","001100100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001000100010","001100100010","010101000100","010101000100","010000110100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001100110011","001000100010"),
		("100110001001","011101100110","001100100010","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001100100010","010101000100","010101000100","010001000100","010000110100","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001"),
		("100110001001","011101100110","001100100010","001000010001","000100010001","001000010001","000100010001","000100010000","001000010001","001000100010","001000100001","001000100010","001100100010","010101000100","010101000100","010001000100","010000110100","001100110011","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000010001"),
		("100110001001","011101010110","001000100010","001000100001","000100010000","000100010001","000100010001","001100100001","010000110010","010100110011","010000110011","001000100010","001100100010","010000110100","010001000100","010001000100","010000110011","001100110011","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001"),
		("100110001001","011101010110","001000100001","001000010001","000100010000","000100010000","001100100010","011101010101","100001010101","100001010101","011000110100","001000100010","001000100010","010000110100","010000110100","010001000100","010000110011","010000110011","001000100010","001000100001","001000100010","001000100010","001000100001","001000100010","001000100001","001000100001","000100010001"),
		("100110001001","011001010110","001000100001","001000010001","000100010001","001000100001","010100110011","011101000100","011000110011","011101000100","100001000101","001100100010","001000100010","010000110100","010000110100","010000110011","010000110011","010000110011","001100100010","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","000100010001"),
		("100110001001","011001010110","001100100010","001100100010","001000100010","001100100010","010000100010","011000110100","011000110011","011101000100","100001010101","001100100010","001000100010","010000110011","010000110011","010000110011","010000110011","010000110011","001100100010","001000100001","001000100001","001000100010","001000100010","001000100010","001100100010","001100100010","001100100010"),
		("100110001001","011101100111","001100100011","001000100010","001100100010","001000100010","001000100001","010100110011","011100110011","011101000100","011101000100","001100100010","001100100010","010000110011","010000110011","010000110100","010000110011","010000110011","001100100010","001000100001","001000100001","001000100010","001000100001","001100100010","011001000100","011101000100","100001000101"),
		("100001111000","100001111000","010101000100","001000100010","001000100010","001000100010","001000100010","010000100010","011000110011","011000110011","010000100010","001000010001","001100100010","010000110011","001100110011","010000110011","010000110011","010000110011","001100100010","001000100001","001000100001","001000100001","001000010001","010000100010","011000110100","011101000101","100001010110"),
		("100001111000","100001111000","011101100110","001100100010","001000100010","001100100010","001100100010","001000010001","001000100001","001000010001","000100010000","000100010000","001100100010","001100110011","001100100010","010000110011","010000110011","001100100010","001000100010","001000100001","001000010001","001000010001","000100010001","001100100010","011000110011","011101000100","100001010101"),
		("100001110111","100001110111","011101100111","010101000100","010001000100","010000110011","001100100010","001000100001","001000010001","001000010001","000100010000","000100010000","001000100001","001100110011","001100100010","001000100010","001000100001","001000100010","001100100010","001100100010","001000010001","000100010000","001000010001","000100010000","001100100010","010100110011","011101000100"),
		("011001100110","011001010110","011101100110","011101100110","011101100111","011101100110","011001010101","010101000100","001000010001","000100010000","000100010000","000100010000","001000010001","001100100010","001000100010","001000100001","001100100010","001100110011","001100110011","001100110011","001000100001","000100010001","001000010001","000100010000","000100010000","001100100010","010100110011"))
	-- 6
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110011010","101010011011","101010101100","101010101100","101010011100","101010101100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100001111001","100001111001","100110001001","101010001001","101010001000","100110001000","101010001010","101010011011","101010101100","101010011100","101010011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001001","100110001010","100101111000","100101010101","100001010100","011000110011","011000110010","011000110011","100001010101","100101111000","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","100001010101","011100110011","011000110010","010100100010","010100100010","010100100010","011000110010","011000110011","100001100111","100110001010","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010101100","101010101100","101010011010","100001010101","010100100010","010000100001","010100100010","010100100010","010100110010","010100110011","010100100010","011101010101","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101110101100","101110101100","101110101100","101010001001","100001000100","011000110011","011000110011","011101000100","100001010101","100001010110","100001010110","011000110011","011001000100","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101100","101110101101","101110101101","100110001001","100001000100","100001010101","100001010101","100001010110","100101100110","100101100110","100101100111","100001000101","011000110100","100110001010","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","100101111000","011101000100","100001010101","100001010101","100001010101","100001010110","100101010110","100101010111","100001010110","011001000100","100110011010","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011010","100001010101","011101000100","011100110100","011101000101","100001010101","011101000101","100001010110","100001010110","011101010101","100110011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110001011","101010011011","101110101100","101110101100","101010011011","100101111000","011101000101","011101000100","011101000100","100001010110","100001010110","100001010110","100101010111","100001010110","100110001001","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110001010","100110011011","101010101100","101110101100","101010011010","100101100111","100001010101","011101000100","011101000101","100001010110","100101100110","100101100111","100101010111","100001010111","100001111001","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001011","100110001010","100101100111","100001010110","011101000100","011101000100","100001010110","100101010111","100101010111","100101010111","100001101000","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110011011","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100101110111","011101000100","011101000100","100001010101","100001010110","100101010110","100101100111","100110001001","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110011011","100010001001","100110001001","100110001010","100110001010","101010011011","101010101100","101010011011","100110001010","100110001010","100110001001","100001010110","100001010110","100001010110","100001010111","100101010111","100101100110","100101111001","101010011010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100110001010","100110011010","101010101100","101010101100","101010011011","100110001001","100001111001","100110001001","100001111000","011001010101","011101010110","100001100110","100001010110","100001010110","100101101000","011101100111","100001111001","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100010001001","100110001001","100001111001","100001111001","100110001010","101010011011","101010101100","101010011011","100101111001","100001111000","100001111000","100001111000","011101100111","011001010101","011101010110","100001010101","100001010110","100001010110","100001100111","010101000100","010000110011","011001010110","100001111000","100110001001","100110001010","100010001001","100001111001"),
		("100110001001","100001111001","100001111001","100001111000","100110001010","101010011011","101010011011","100110001010","100001111000","100110001001","100110001010","100001111001","100001100111","011001000101","011101010110","100001010101","100001010110","100001010110","100001111000","010101000100","001100100010","001100100010","001100100010","010000110011","010101000100","011001010110","011101100111"),
		("101010011011","100110001010","100001111001","100001111001","100010001001","100110011010","100110001010","100001111000","100001111001","100110001010","100110001010","100110001001","011101100110","010101000101","011001010101","011101010101","100001000101","100001010110","100110001001","010101000100","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010"),
		("101010011011","100110001010","100001111001","100010001001","100010001001","100001111001","100001111001","100001111000","100010001001","100110001010","100101111001","011101100110","100001100111","011001010110","011001010101","011101000101","011101000101","100001111000","100001111001","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","100001100111","010100110011","010100110011","100001111000","100001111000","011101010101","011101000100","100001100111","100110001010","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111000","100001111001","100110001001","100110001010","100001111001","100110001001","011101010110","010000110011","001100100010","001100100010","100001100111","100001111000","011101100111","011101010110","100001100111","011101111000","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001001","100001111001","100010001001","100110001010","101010011010","100101111000","011001000101","010000100010","001000100010","001000100010","001000100010","011001010101","100001111000","011001010110","011001010101","011001010101","010101000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100110001001","100110001010","100101111000","010100110011","001100100010","001100100010","001000100010","001000100010","001000100001","001100100010","011101100110","011001010110","010101010101","010101010101","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100110001001","100110001001","011101100111","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","010001000100","010101000101","011001010101","010101000101","001100110011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010"),
		("101010011011","100110001001","100010001001","100110001001","100110001001","011101100110","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101000101","010101010101","010101000100","001100100011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100110001001","101010011010","011101100111","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010001000100","010101000101","010101000101","010101000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","101010011010","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","010001000100","010101000100","010101000101","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001"),
		("100110001001","100010001001","100110001001","100110001001","100110001001","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110100","010001000100","010101000101","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100010001001","100010001001","100010001001","100110001001","100001111001","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","010000110011","010101000100","010000110100","010000110011","010100110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001001","100110001001","100110001001","100110001001","100110001010","100001111001","001100100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","010000110011","001100110011","010000110100","010000110011","010100110100","100001000101","011101000100","010100110011","001100100010","001000100010","001000100010","001000100001","001000010001","001000100001"),
		("100110001010","100010001001","100110001001","100110001001","100110001010","100110001001","010000110010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","001100100010","010000110011","010000110011","011101000101","100001010101","100001010101","100001010101","010100110011","001000100010","001000100010","001000100001","001000010001","001000010001"),
		("100110001001","100110001001","100010001001","100110001001","100110001010","100110001010","010000110011","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","010000110011","001100100010","010000110011","010000110011","011001000100","011101000100","100001010101","100001010101","100001000101","010000100010","001000100001","001000100001","001000100001","001000010001"),
		("100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","010101000100","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","010000110011","001100100010","010000110011","010000110011","010100110011","011101000100","100001000101","100001010101","100001010101","011001000100","001000100001","001000100010","001100110011","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","100110001001","100101111001","010101000100","001000100001","001000010001","001000100001","001000100001","001000100010","001000100001","010000110011","001100100010","010000110011","010000110011","010000110011","011000110011","100001000101","100001010101","100001010101","011001000100","001000100010","001000100010","001100100010","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","100110001001","100101111000","011001000101","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","001100100010","010000110011","010000110011","001100100010","010000100010","011000110011","011101000100","100001000101","011001000100","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100110001001","100101111000","100101111000","100001100111","010101000100","001100100010","001000100001","001000010001","001000010001","001000100001","001000100001","010000110011","001000100010","001100110011","001100100010","001000100010","001000100001","001000100001","001100100001","010000100010","001100100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100101111001","100001100111","100001000101","011101000100","010100110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","010000110011","001000100010","001100100010","001100100011","001100100010","001000100010","001000100001","001000010001","000100010000","001000010001","001000100010","001100100010","001000100010","001000100010"),
		("100110001001","100001110111","100001010101","100001010110","011101000101","010100110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","001000100001","001000100010","001100100010","001100100010","001000100001","001000100001","001000010001","000100010000","001000010001","001100100010","001100100010","001000100001","001000100001"),
		("100110001001","100001111000","011101000101","100001010110","100001010101","011000110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000010001","000100010000","000100010001","001000010001","001000010001","001000010001","001000010001"),
		("100010001001","100001111000","011101010110","011101000101","100001000101","011000110011","001000100001","000100010001","000100010000","000100010001","001000010001","001000010001","001000100001","001100110011","001100100010","010000110100","010001000100","010001000100","010000110011","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100010"),
		("100001111000","100001111000","011101010110","011000110011","011000110011","001100100010","001000100001","001100110011","010101000101","001100110011","000100010000","001000010001","001000010001","001100110011","001100100010","010101000100","010101010101","010101010101","010101000100","001000100001","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","011101100110","010000110011","010000110011","010101000101","011101100110","100001111000","100001111000","010001000100","001000010001","000100010000","001000010001","001100110011","001100100010","010101000101","010101000101","010101010101","010101000100","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100001110111","100001110111","100001100111","011101100111","100001111000","100001111000","100001111000","100001111000","011001010110","010101000100","001000010001","000100010000","001000010001","001100100010","001100100010","010101000101","010101000101","010101000101","010101000100","001100100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("011001100110","011001100110","011101100110","011101100110","011101100111","011101100110","011101100111","011001010110","010000110011","001000100001","000100010000","000100010000","001000010001","001100100010","001100100010","010101000100","010101000100","010101000100","010101000100","001100100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"))
	-- 7
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100010001001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100101100110","100001010101","100001010100","011101000011","011101000100","100001100111","100110001001","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111001","100001100111","011100110011","011000110010","010100100010","010100100010","010100100010","011000110010","011101000100","100101111001","100010001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100101111001","100101010101","011000110010","010000100001","010000100001","010100100010","010000100001","010100100010","010100100010","011101000101","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100101111000","100001010100","011000110011","011000110011","011000110011","011000110011","011001000100","011000110100","010100100010","011000110011","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100001111001","100001111001","100101100110","100001000100","100001000101","100001010101","100001010110","100101100110","100101100111","100101100111","011001000100","011000110100","100110001010","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001001","100110001010","100110001001","100001010101","011101000100","100001010101","100001010101","100001010110","100101100110","100101100111","100101100111","011101000101","011000110100","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","101010011011","100101100111","100001000101","011101000100","011101000100","100001010101","100001010101","100001010101","100001010110","011101000101","011101000101","100110001010","100010001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010101100","101010101100","101010101100","101010011100","100110001001","100001100110","011101000100","011101000100","011101000101","100001010110","011101000101","100001010110","100001010101","100001100111","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101110101100","101110101100","101110101100","101010011100","101010011011","100101100111","100101100111","011101000101","011101000100","011101000101","100101010110","100101100110","100101100111","100001010110","100001100111","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101100","101110101101","101110101100","101010011011","101010011011","100101101000","100001100110","011101000101","011101000100","011101000101","100001010110","100101100111","100101010111","100101010110","100101111000","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","101010011011","100110001010","100101111000","100001010101","011101000100","100001000101","100101010110","100101010111","100101010111","100101101000","100110011010","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","101010011011","101010011011","100110001001","100001010101","011101000100","011101000100","100001010110","100001010110","100101010110","100110001010","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110001011","101010011011","101110101100","101110101100","101010101100","101010011011","100110001010","100001111001","100001100110","100001000101","100001010101","100101100110","100101010111","100001010110","100110001001","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110001010","100110011011","101010101100","101110101100","101010011011","100110001010","100001111001","100001111001","100001100110","011101000100","011101000100","100001000101","100101010110","100101010111","011101100110","011101100111","101010011010","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100001111001","100110001001","100001100111","011101000100","011101000100","100001010110","100101010111","100101100111","011001010110","001100100010","011001010101","100001111000","100001111000","100001111001","100110001010","100010001001"),
		("101010101100","101010011011","100110001010","100110001010","100110011011","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100110001010","100110001010","100001010101","011101000100","011101000100","100001000101","100001010110","100101111001","011001010110","001100100010","001100100010","010000110011","010000110011","011001000100","011001010101","011001010110"),
		("101010011011","100110011011","100010001001","100110001001","100110001001","100110001010","101010011011","101010101100","101010011011","100110001010","100110001001","100110001001","100101111001","100001010110","100001010110","100001010101","011101000100","100001100111","100110001010","010101000101","001100100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100110001010","100110001010","100110011010","101010101100","101010101100","101010011011","100110001001","011101100110","011101010101","100101111000","100001100111","011001010101","011101010101","100001010110","100110001001","100001111000","001100110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010101100","101010011010","100001111000","011001000100","010000100010","010100110011","100101111000","011101100111","011001000101","011101100110","100001111001","100110001010","010101000101","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100001111001","100001111001","100001111000","100110001010","101010011011","101010011010","100001100111","010100110011","001100100010","001100100010","010000110010","100001100111","011101010110","011001010101","011001010110","011001010110","011001010101","001100100011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111001","100010001001","100110001010","011001010101","010000100010","001100100010","001000100010","001000100010","001000100010","010000110011","011001010101","011001010101","011001010110","011001010101","010001000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100010001001","100110001001","100001111000","010000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","011001010101","011001010101","010101010101","010000110011","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100010001001","100001111001","100001111001","100001111000","010000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","011101100111","011001010101","010101000101","001100110011","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111001","100110001001","100001111000","010000100010","001000100010","001000100001","001000100010","001100100010","001100100010","001000100010","010101000101","100001100111","011001010101","010101000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001001","100001111001","100010001001","100110001010","100110001001","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000101","100001111000","010101000101","010001000100","001100100010","001100100010","001100100011","001100100010","001100100010","001100100010","001000100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100110001001","100110001010","100110001010","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","011001010110","010101000100","010000110011","011001000100","100001010101","100001010101","011101000101","010100110011","001000100010","001000100010","001000100010","001100100010","001000100010"),
		("101010011011","100110001010","100010001001","100110001001","100110001001","100110001010","010100110100","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","010000110011","010101000101","010001000100","001100100010","011001000100","100001000101","100001000101","100001000101","100001000101","010000110011","001000100010","001000100010","001100100010","001000100010"),
		("101010011011","100110001001","100010001001","100110001001","100110001001","100101111001","010100110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101000101","010000110100","001100100010","010000110011","011101000101","100001000101","100001000101","100001010110","100001000101","001100100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100110001001","101010011010","100101111001","010101000100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101000100","010000110011","001100100010","001100100010","011100110100","011101000100","100001000101","100001010110","100001010110","010000110011","001000100001","001000100010","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","100110011010","100101111000","011001000101","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","010000110100","010101000100","010000110011","001000100010","001000100010","001100100010","010000100010","010100110011","011101000101","100001010110","010100110011","001000100001","001000100001","001000100001"),
		("100110001001","100010001001","100110001001","100110001001","100001111001","100101111000","100001100111","001100100011","001000100010","001000100010","001000100010","001000100010","001000100010","010000110100","010101000100","010000110011","001000100001","001000100001","000100010001","000100010000","000100010000","010000100010","010100110011","010000100010","001000100010","001000100001","001000100001"),
		("100110001001","100110001010","100010001001","100110001001","100001111000","100110001001","100110001001","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","010101000100","001100110011","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010001","000100010001","001000100001","010000110011","010001000100"),
		("100110001010","100110001010","100110001001","100110001001","100110001001","101010011011","100110001010","010001000100","001000100001","001000100001","001100110011","001000100010","001000100001","010000110011","010101000100","001100100010","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001000010001","001100100010","001100110010"),
		("100110001010","100110001001","100110001001","100110001001","100110001001","101010011010","100101111001","010000110011","001000100010","001100100010","010000110100","001000100010","001000100010","010000110011","010101000100","001100100010","001000100001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001"),
		("100110001001","100110001001","100010001001","100110001001","100110001010","101010011010","011101100111","001100100010","001000100001","001100100010","010000110011","001000100010","001000100010","010000110011","010000110011","001000100010","001000010001","001000010001","001000010001","001000010001","000100010000","001000100001","001100100010","001000010001","001000010001","001000010001","001000010001"),
		("100110001001","100110001001","100110001001","100110001001","100001100111","100001010110","010100110011","001000100001","001000100001","001000100001","001100100010","001000100001","001000100001","001100100011","010000110011","001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000100001","001000010001","000100010001","001100110010","001000100001"),
		("100110001001","100110001001","100010001001","100001100111","100001000101","011101000100","010100110011","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001100110011","010000110011","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010"),
		("100110001001","100110001001","100001111000","100001010110","100001010110","100001010101","011000110011","001000100001","001000010001","001000010001","001000100001","001000010001","001000010001","010000110011","001100110011","001000010001","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100110001001","100101111000","100001010110","100001010110","100001010110","011000110100","001000010001","001000010001","001000100010","001000100001","001000100001","001100100010","010101000100","010000110011","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001001","100110001001","100001100111","100001000101","100001000101","011000110011","010001000100","011101100111","011001010101","001000010001","001000010001","001100100010","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100010001001","100001111000","011101000101","011101000101","011101100111","100001111001","100110001001","010001000100","000100010001","001000010001","001100110010","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001001","100010001001","100010001001","100010001001","100110001001","100001111001","100001111000","100001111000","100001111000","001100100010","000100010001","001000010001","001100110011","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100010001001","100001111001","100001111000","100001111001","100110001001","100001111000","100001111000","100001111001","011101100111","001000100010","000100010001","001000010001","010000110011","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100110001001","100110001001","011001010110","001000100001","001000010001","001000010001","010000110011","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","100001110111","100001111000","100001111000","100001111000","100001111001","100001111001","010000110100","001000100001","001000010001","001000010001","010000110100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100001110111","100001100111","100001100111","100001100111","100001111000","100001111000","100001111000","011101100111","010000110011","001000100001","001000010001","001000010001","010100110100","010101000100","010000110011","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100001","001000100010","001000100010"),
		("011001100110","011001100110","011101100110","011101100110","011101100111","011101100110","011101100111","010101010101","001100100010","001000010001","000100010000","001000100001","010000110100","010000110011","010000110011","001000100010","001000100001","001000010001","001000100001","001000100001","001000100001","001000100010","001000100001","001000100010","001000100001","001000100010","001000100010"))
	-- 8
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100010001001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100001111000","100101010101","100001010100","011101000100","011101000100","011101010101","100001111000","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111001","100001111000","100101100110","011000110010","010100100010","010100100010","010100100010","010100100010","011000110011","100001100111","100010001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100001111001","100101100111","100001000100","010100100010","010000100001","010000100010","010000100001","010000100010","010100100010","011000110011","100101111000","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110001001","100101100110","100001000100","011000110011","011000110011","011000110011","011000110011","011000110011","010100110010","010100100010","100001111000","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100001111001","100001111001","100101111000","011101000100","100001010101","100001010101","100001010110","100101010110","100101100111","100101100110","100001010101","010100100010","100001111000","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001001","100110001010","100110001001","100001100111","011101000100","100001010101","100001010101","100001010110","100101100110","100101100111","100101100111","100001010110","011000110011","100001100111","100010001010","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","101010011011","100101111000","100001010101","100001010101","011100110100","011101000100","100001010101","100001010110","100001010110","100001010110","011000110100","100001111001","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010101100","101010101100","101010101100","101010011011","100101111000","100101100111","011101000101","011101000100","011101000100","100001010110","011101000101","011101000101","100001010101","011101010110","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101110101100","101110101100","101110101100","101010101100","101010011011","100001010110","100101100110","100001000101","011101000100","011101000100","100001010110","100101100110","100101100110","100001010110","100001101000","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101100","101110101101","101110101100","101010011011","101010011011","100101111000","100101100110","011101000101","011101000100","011101000100","100001010110","100101010110","100101010111","100101010110","100101111000","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","101010011011","101010011010","100101111000","100001010101","011101000100","100001000101","100001010110","100101010111","100101010111","100101100111","100110001010","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","101010011011","101010011011","100110001001","100001010101","011101000100","011101000100","100001010110","100001010110","100101100111","100110001010","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110001011","101010011011","101110101100","101110101100","101010101100","101010011011","100110001010","100001111000","100001010101","011101000101","100001010101","100101010110","100101010110","100101100111","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110001010","100110011011","101010101100","101110101100","101010011011","100110001010","100001111001","100001100111","011101000100","011101000100","011101000100","100001010101","100101010110","100101100111","100001111001","100110001010","101010011010","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100001111001","100001100110","100001000101","011101000100","100001010101","100001010110","100101010111","100001100111","011001010101","100110001001","101010011010","100110001010","100001111001","100001111001","100110001001","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110011011","100110001010","100110001010","100110001010","100110001001","100001111001","100010001001","100101111000","100001000101","011101000100","011101000100","100001000101","100001010101","100101100111","011101100110","001100100010","010001000100","011101100110","100001100111","100001111000","100001111001","100110001001","100001111001"),
		("101010011011","100110011011","100010001001","100110001001","100110001010","100110001010","101010011011","101010011011","100001111000","011101010110","100001100111","100101111000","100001010110","100001010110","011101000101","011101000101","100001010110","100110001001","011001010110","001100100010","001100100010","001100100010","010000110011","010101000100","011001010101","100001100111","100001111000"),
		("101010011011","100110001010","100010001001","100110001010","100110001010","100110001010","100101111000","011101010101","010100110011","010100100010","100001010110","100101111000","011001010101","011001010101","011101010101","100001100110","100110001001","100010001001","010000110100","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","010000110011"),
		("100110001010","100110001010","100001111001","100010001001","100001100111","011001000101","010100110011","001100100010","001100100010","001100100010","100001010110","100101111000","011001010101","011001010101","100001110111","100110001010","100110001010","011001010110","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100001111001","100001111001","100001111001","010101000100","001100100010","001100100010","001000100010","001100100010","001100100010","010000110011","010101000100","011001010101","011001010101","011101010110","011101100111","100001111000","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111000","010000110011","001100100010","001000100010","001100100010","001100100010","001000100010","001000100001","010000110011","011001010101","011001010101","011001010101","011001010101","010101000101","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100001111000","010000110011","001000100010","001100100010","001100100010","001000100010","001000100010","001000100001","010000110011","011001010101","011001010101","011001010101","011001010101","010001000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111000","010000110011","001000100001","001100100010","001000100010","001000100010","001000100010","001000100001","010000110011","011001010110","011101100110","011001010101","010101000101","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111000","010000110011","001000100001","001100100010","001000100010","001000100001","001000100010","001100100010","010000110011","011101100110","011101100111","010101010101","010101000100","001100100011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001001","100001111001","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","011101100111","011101100111","010101000101","010101000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001010","100110001001","011101100110","001100100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100001","001100110011","011001010110","011001010101","010101000100","010000110100","001000100010","001000100010","001000100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001"),
		("101010011011","100110001010","100110001001","011101100110","001100100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100001","001100100010","010101000100","010101000100","010101000100","010000110011","001000100010","001000100010","001100100010","011101000100","011101000101","011001000100","010100110011","001100100010","001000100010","001000100010","001000010001"),
		("101010011011","100110001001","100001111001","011101100110","001100100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","010101000100","010001000100","001100100010","001000100010","001000100010","001100100010","011100110100","100001000100","100001010110","100001010110","011001000100","001000100010","001000100010","001000010001"),
		("100110001010","100110001001","100110001001","011101100111","001100100010","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","010101000100","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","010100110011","011101000100","100001010110","100001010110","100001010101","010000110011","001000100001","001000100001"),
		("100110001001","100110001001","100110001001","011101100110","001100100010","001000100001","001000010001","001000100001","001000100010","001000100010","001000100001","001000100001","010000110100","010101000100","010000110011","001100100010","001000100001","001000100010","001000100001","001100100010","011100110100","100001000101","100001010110","100001010110","011001000100","001000100001","001000100001"),
		("100110001001","100010001001","100110001001","011101010110","001100100010","001000100001","001000100001","001000010001","001000100010","001000100010","001000100010","001000100010","010000110011","010101000100","010000110011","001000100010","001000100001","001000100001","001000010001","001000010001","010000100010","011000110100","011101000101","100001010101","011101000101","001100100010","001000100001"),
		("100110001001","100110001010","100110001001","011001010110","001100100010","001000100001","001000100001","001000010001","001000100001","001000100010","001100100010","001100100010","010000110011","010101000100","010000110011","001000100001","001000100001","001000100001","001000010001","000100010001","000100010001","000100010000","001100100001","011101000100","011101000100","001100100010","001000100010"),
		("100110001010","100110001010","100110001001","011101010110","010000110011","001100100010","001100100010","010101000100","011101010101","011101000100","011100110100","010100110011","010000110011","010101000100","001100110011","001000100001","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010000","001000010001","001000100001","001000010001","001000100001"),
		("100110001010","100110001001","100110001001","100001111000","010000110011","001100100010","010101000100","100001010110","011101000100","011100110011","011100110011","010100100010","010000110011","010101000100","001100110011","001000100001","001000100001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001"),
		("100110001001","100110001001","100110001001","100010001001","010100110011","010000100010","001100100010","010100110100","011101000100","011100110011","011100110011","010100100010","010000110011","010101000100","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","000100010001","001000010001","001000010001","001000010001","001000010001"),
		("100110001001","100110001001","100110001001","100110001001","011101010110","001100100010","001000100010","010000100010","011100110011","011000110011","011000110011","010000100010","010000110011","010001000100","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","001100110010","001000100001"),
		("100110001001","100110001001","100110001001","100110001001","100001111001","011101010110","010100110100","001100100001","010100110011","011000110011","010100100010","001000010001","010000110011","010000110100","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001"),
		("100110001001","100110001001","100110001001","100110001001","100110001010","100101111001","100001100111","010100110011","001100100001","001000100001","001000100001","001000010001","001100110011","010000110011","001000100010","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","101010011010","100110001010","100101111000","100001111000","011001010110","001100110011","001000010001","001000010001","001100100010","001100100010","001000010001","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100110001001","101010011010","101010011010","100110001001","100001111000","011101100111","010000110011","001000010001","001000100010","010000110011","010000110011","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100010001001","100110001001","101010011010","101010011010","100001111001","100001111000","011101100111","001100110011","001000100001","010000110011","010101000100","010000110100","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001001","100010001001","100010001001","100010001001","101010011010","100110001001","100001111000","100001111000","011001010101","001100100010","001000100001","010000110100","010101000100","010101000100","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100010001001","100001111001","100001111000","100001111001","100110001001","100001111000","100001111000","100001111000","010101000100","001000100010","001000100010","010101000100","010101010101","010101000100","001000100010","001000100001","001000010001","001000010001","001000010001","001000100001","001100100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100110001001","011101100111","001100110011","001000100001","001000100010","010101000101","010101010101","010101000101","001100100010","001000100001","001000010001","001000010001","001000010001","001000100001","001100110011","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","100001110111","100001111000","100001111000","100001111000","100010001001","011001010110","001100100010","001000100001","001100100010","010101010101","010101010101","010101010101","001100110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001110111","100001100111","100001100111","100001100111","100001111000","100001111000","100001111000","011001010101","001100100010","001000100001","001000100010","010101010101","010101000101","011001010101","010001000100","001000100001","001000010001","001000010001","000100010000","000100010001","000100010001","001000010001","001000010001","001000100010","001000100001","001000100010","001000100010"),
		("011001100110","011001100110","011101100110","011101100110","011101100111","011101100110","011101100111","010101000100","001000100010","001000010001","001000100001","010101000101","010101000100","010101000101","010101000100","001000100001","001000010001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100001","001000100010","001000100010"))
	-- 9
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","100110011010","100110001010","100110001001","100010001001","100010001001","100010001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111001","100001110111","100101100110","100101100110","100001100110","100101110111","100110001001","100110001001","100110001001","100110001010","100010001001","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100101111000","011101000011","011000110010","011000110010","010100100010","010100100010","011000110011","100001100111","100110001001","100101111001","100110001001","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100101100101","011000110010","010000100001","010000100001","010100100010","010100100010","010100100010","011100110011","100101111000","100110001001","100110011010","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100010001001","100101110111","100001010100","011000110010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","100001010110","100110001001","100110001010","100110011010","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001010","100110001010","100001100110","011101000011","100001000100","100001010101","100001010101","100001010101","100001010110","100001010101","010100110011","011101010101","100010001001","100001111001","100001111001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","011101000101","011101000011","100001010101","100001010101","100101100110","100101100110","100101100110","100101100111","011101000100","011101010110","100110001010","100110001010","100010001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010101100","101010101100","101010011011","100001010110","011101000100","011101000100","011101000100","100001010101","100101010110","100101010110","100101100111","011101000100","100001100110","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101110101100","101110101100","101110101100","101010011011","100101100111","100001000101","011101000100","011101000100","011101000101","100001010101","011101000101","100001010110","011101000101","100101111001","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101100","101110101101","101110101100","100101111000","100001010110","100101100110","100001000101","011101000101","100001000101","100101010110","100001010110","100101010110","100001100110","101010011010","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","100110001001","100001010101","100001010110","100001000101","011101000101","011101000100","100001010110","100101100111","100101010110","100001100111","100110001010","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","100101111001","100001010110","011101000100","011101000100","100001010101","100101010110","100101010110","100001010110","100101111000","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110001011","101010011011","101110101100","101110101100","101010101100","101010011011","100001010110","011101000100","011101000100","011101000101","100001010110","100101010110","100101100111","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110001010","100110011011","101010101100","101010101100","101010011011","100110001010","100001010110","011101000101","011101000101","100001010101","100101100110","100001010110","100001111000","100001111000","100001111000","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100001111000","100001000101","011101000100","011101000100","100001000101","100001010110","100001010110","100101111000","100001111000","100001111000","100110001001","100110001010","100110001010","100001111001","100001111001","100110001001","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110011011","100110001010","100110001010","100110001010","100010001001","100001111001","100001111000","100001000101","011101000100","011101000100","100001010101","100001010110","100001010110","100001111000","100110001001","100110001001","100001111001","100001111000","100001111000","100001111000","100001111001","100110001001","100001111001"),
		("101010011011","100110011011","100010001001","100110001001","100110001001","100110001010","101010011011","101010011011","100110001001","100101111000","100001100110","011101000101","100001010110","100001100110","100001010110","100001010110","100101100111","011001010101","011001010110","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000","100001111000"),
		("101010011011","100110001010","100010001001","100110001010","100110001010","100110001001","100101111000","011101010110","011101000101","100001100111","100001100110","011101000100","011001010101","011001010101","011101010101","100001010110","100101111001","010101000101","001100100010","010000110100","011001010110","100101111000","100110001010","100110001010","100110001001","100001111000","100001111000"),
		("100110001010","100110001010","100001111001","100001111000","100001100111","011001000101","010100110011","001100100010","001100100010","100001100111","100101111000","011101010101","011001010101","011001010101","011101100110","100001111000","100110001010","010101000100","001100100010","001100100010","001100100010","001100110011","010101000101","100001100111","100110001001","100010001001","100001111000"),
		("100110001010","100001111001","011101100110","011001000100","010000110011","001100100010","001100100010","001000100010","001100100010","100001100111","100110001001","100001111000","010101010101","011001000101","100001111000","100110001010","011101100111","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001100100010","010101000100","100001110111","100001111001"),
		("101010011011","100001111001","010000110011","001100100010","001100100010","001100100010","001000100010","001100100010","001100100010","011101010110","011101100111","011101100111","010101010101","010101010101","100001111000","100001111001","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","011101100111"),
		("101010011011","100001111000","001100100010","001000100010","001100100010","001000100010","001100100010","001100100010","001000100010","001000100010","010001000100","011001000101","011001010101","011001010101","011101100111","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100"),
		("101010011011","011101100111","001100100010","001000100010","001100100010","001000100010","001100100010","001000100010","001000100010","001000100010","010001000100","010101000101","011101010110","011101100110","011001010110","010001000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","010000110011"),
		("101010011011","011101100110","001100100010","001000100010","001100100010","001000100010","001100100010","001000100010","001000100001","001000100010","010101000100","010101000101","011101100110","011101100111","011001010101","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100011"),
		("101010011011","011001010101","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101000101","011101100111","011101100111","010101000101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001100100010","001100100010","001100100010"),
		("101010011011","010101000100","001000100001","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","010000110100","010101000101","011001010101","011001010110","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","010101000100","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","010000110011","011001010101","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","010001000100","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","010000110011","010101000101","010101000100","010101000101","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","010000110100","001000100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100010","001000100010","001100110011","010101000101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100001","001100100010","010000110011","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","010000110011","001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001000100010","001000100010","001100100010","010101000100","010101000100","010001000100","001000100010","001000100010","001000100010","001000100010","001000100001","010000100010","011101000100","011000110011","010000100011","001000100010","001000100010","001000100001","001000100001"),
		("100001100111","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000100010","001000100010","001100100010","010101000100","010101000100","010000110011","001000100001","001000100001","001000100001","001000100001","001000100010","010100110011","011101000100","100001000101","100001010101","010000110011","001000100001","001000100001","001000100001"),
		("011101100110","001100100010","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010000110100","010101000100","010000110011","001000100001","001000100001","001000100001","001000100001","001000010001","010100110011","011101000100","100001000101","100001010110","011000110100","001000100001","001000100001","001000100010"),
		("100001100111","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010101000100","001100110011","001000100001","001000100001","001000100001","001000010001","001000010001","010000100010","011100110100","011101000101","100001010110","011000110100","001000100001","001000100001","001000100001"),
		("100001100111","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010101000100","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","010100110011","011101000101","100001010101","010000110011","001000100001","001000010001","001000100001"),
		("100001111000","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110100","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","000100010001","001100100001","011000110011","011000110100","001100100010","001000100001","001000100001","001000100001"),
		("100101111001","011101010110","001100100010","001000100001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","010000110011","010000110100","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100001","001100100001","001000100001","001000100010","001100110011","001000100010"),
		("100110001001","011101010110","001100100010","001100100010","010000110011","010100110011","010100110011","010000110010","001000100001","001000010001","001000010001","001100110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010"),
		("100110001001","011101010110","001000100001","010000110011","011101010101","100101100110","100001010101","011101000100","001100100001","001000100001","001000100001","001100100010","010000110011","001100100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010"),
		("100110001001","100001111000","010000110011","010000110011","100001010101","100001000101","011101000100","011000110011","001100100001","001000010001","001000010001","001000100010","001100110011","001100100010","001000010001","001000100001","001000010001","001000010001","001000100001","001000100010","001000010001","000100010001","000100010001","001000010001","001000100001","001000100001","001100110011"),
		("100110001001","100110001001","100001111000","010101000100","011000110100","011000110011","011000110011","011000110011","001100100001","000100010001","001000010001","001000010001","001100100010","001100100010","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","000100010000","001000010001","001100110011","010000110011","010101000101","100001111000"),
		("100110001001","100010001001","100110001001","100001111000","011101000101","011000110011","011100110011","011000110011","001000100001","001000010001","001000010001","001000010001","001100110010","001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010001","001100100010","100001110111","100110001001","100110001001","100110001001"),
		("100110001001","100010001001","100010001001","100010001001","100001111000","011000110011","011000110011","010000100010","001000010001","001000010001","001000010001","001000100010","001100110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001100100010","011101100111","100110001001","100110001001","100110001001"),
		("100010001001","100001111000","100001111000","100010001001","011101100111","001100100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000100001","001100110010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","010101000101","100110001001","100110001001","100110001001"),
		("100001111000","100001111000","100001111000","100001111000","010101000101","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001100110010","001000100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100001","010000110100","100001111001","100110001001","100110001001"),
		("100001111000","100001111000","100001111000","100001111000","010000110011","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001100110011","001100100010","001000010001","001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","001000100001","001000010001","010000110011","100001111000","100010001001","100010001001"),
		("100001110111","100001100111","100001110111","011101100111","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","001100100010","001000100010","001000010001","001000010001","001000010001","001000010001","001100110011","001000100001","000100010001","001000010001","001000010001","001100100010","011101100111","100001111000","100001111000"),
		("011001100110","011001100110","011101100110","011001010101","001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001100100010","011001010110","011101100111","011101100111"))
	-- 10
	,

		(	("101010011100","101010101100","101010101100","101010101100","101010101100","100110011011","100101110111","100101100101","100101100101","100001010100","011100110011","010000100001","010000100001","010000100001","010000100010","001100100001","001100010001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","010000100010"),
		("101110101100","101110101101","101110101100","101110101101","101010101100","100101111000","100101010101","011101000011","011101000011","011100110011","010100100010","001100100001","001100010001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","010000100001","010000100010"),
		("101110101100","101110101100","101110101100","101110101100","101010001001","100101100101","011101000011","010100100010","010100100010","010100100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100001","010000100010","010000100010","010000100010","010000100010","010000100001","001100100001","010000100010","010000100001"),
		("101110101101","101110101101","101110101101","101110101100","100101100110","100001010100","100001000011","011000110011","010100100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","010000100001","010000100010","010000100010","010100100010","010000100010","010000100001","010000100001","001100100001","001100100001","010000100001","001100100001"),
		("101010101100","101010011100","101010011011","100110001010","100101010101","011101000011","011101000011","010100110010","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100100001","010000100001","010000100010","001100100001","010000100001","010000100001","010000100001","001100100001","001100010001","001100100001","001100100001","001100100001"),
		("100110001010","100110001011","100110011011","100101111001","100101100110","011101000011","010100100010","010000100001","010000100001","010000100001","010000100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001"),
		("100110001011","100110011011","100110011011","100110001010","100101111001","100001100110","010100100010","010000100001","001100100001","010000100001","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100101100111","011100110011","010100100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100001","010000100010","001100100001","001100100001"),
		("100110011011","100110011011","100110011011","100110001010","100110001011","100110001001","100001000101","011000110010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100010","010000100010","010000100010","010100100010","010000100010","010000100010","010000100010","010000100010"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","100110001010","100101111000","011101000100","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010100100010","010100110011","010100110011","011000110011","011000110011","010100110011","010100110011","010100100010"),
		("100110011011","100110011011","100110011011","100110011011","100110001010","100110001010","100110001001","100101100111","011000110011","010100100010","010000100001","010000100001","001100100001","010000100001","010000100001","010000100010","010000100010","010100100010","011000110011","011000110100","011101000100","011101000101","011101000101","011101000101","011101000100","011000110011","010100110011"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100110001010","100101111001","011101000101","011000110011","010100110011","010000100010","010000100010","010100100010","010100110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010101","100001010101","100001010110","100001010110","100001000101","011101000100","011000110011"),
		("100110001010","101010011011","101010011011","100110011011","100110001010","100001111001","100010001001","100101111001","100001010101","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110100","011000110100","011101000100","100001000101","100001010101","100001010110","100001010110","100001010110","100001010110","100001010110","011101000101","011000110011"),
		("101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001","100001111000","011101000101","011101000100","011101000100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","011101000101","011000110011"),
		("101010101100","101010101100","101010011100","101010011011","100010001001","100001111001","100001111001","100001100111","011101000100","011101000100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100101010111","011101000101","011000110100"),
		("101010101100","101110101100","101010101100","101010011011","100010001001","100001111001","100001111001","100001100111","011101000100","011101000100","011000110100","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110","100101010111","100001010101","011101000100"),
		("101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","100010001010","100001100111","011101000100","011001000100","011000110100","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001010110","100001010110","100001010111","100001010110","011101000100"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","100110001011","100110001010","100101100111","100001000101","011101000100","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010111","100001010110","011101000100"),
		("101010011011","101010011011","101010011011","101010011011","100110011011","100110011010","100110001001","100101100111","100001010101","011100110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010111","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100101100111","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110","100001010111","100001010111"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","100110011011","100110001001","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000101","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101010101100","101010011100","100110001001","100001100110","011000110011","010100100010","010100110010","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","101110101100","100110001010","100101111000","011101000101","011000100011","010100100010","010100100010","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000101","100001010110","100001010110","100001010111"),
		("101110111101","101110111101","101110111101","101110101101","101110111101","101010101100","100110001010","100010001001","100001010110","011000110011","010100100010","010100100010","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","011000110011","011101000100","100001000101","100001010110","100001010111"),
		("101110111101","101110111101","101110111101","101110101101","101110101101","101010011100","100110001010","100010001001","100101100111","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000100","100001000101","100001010110","100101010111"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010101100","100110001010","100110001001","100101100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","011000110011","011000110100","011101000100","011101000100","100001000101","100001010110","100101010111"),
		("101110101101","101110101101","101110101101","101110101101","101110111101","101010011011","100110001010","100110001001","100001010110","011000110100","011100110100","011100110100","011101000100","011101000100","011101000100","011000110011","011000110011","011000110011","011000110010","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110","100001010111"),
		("101110111101","101110101101","101110101101","101110101101","101110101101","101010011011","100110001010","100110001001","100001010101","011000110100","011101000100","011101000100","100001010110","100001010110","100001000101","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010011100","100110001010","100110001001","100001010110","011101000100","100001010101","011101000101","100001010110","100001010111","100001010110","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101110111101","101010011011","100110001010","100110001010","100001100111","100001010101","011101000101","011101000101","100001010110","100001010111","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100110001010","100101111000","011101000101","011000110100","011101000101","100001000101","100001000101","100001010110","011101000100","011000110010","010100100010","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","100110001001","011101000100","011000110011","011100110100","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010011010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001010101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","101010011011","101010011011","011101010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010101","100001010110","100001010110","100001010110"),
		("101110111101","101110111110","101110111110","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","100001111000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010101","100001010101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011100","101110101101","101010011010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001010101","100001010110","100001010110"),
		("101110111101","101110101101","101110101101","101110101100","101010011011","100110011011","100110011011","101010011011","101010101100","101010101100","100001101000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110010","011000110011","011000110011","011100110100","100001000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111101","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","101010101100","101110101100","101110101100","101010011011","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001010101","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","100110011011","100110011011","100110011011","101010101100","101010101100","101010101100","101010101100","100101111000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","100001000101","100001010101"),
		("101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","100110011011","101010101100","101110101100","101010101100","101010011100","100110001010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","011101000100","011101000100","011101000101","100001000101","100001000101"),
		("101110111101","101110111101","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","101110101101","100001111001","010100110100","010101000100","010101000100","010101000100","010101000100","011001000100","011101100110","011101000101","011000110011","011000110100","011101000100","100001000101","100001000101","100001000101","100001000101","100001000101","100001000101"),
		("101110111101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011011","101110101101","101110101101","011101100111","010000110011","010000110011","010001000100","010101000100","010101000101","010101000101","011101100111","011101010110","011000110100","011101000100","011101000100","011101000101","011101000101","011101000100","011101000100","011101000100","011101010101"),
		("101110101101","101110111101","101110111101","101010011011","100110011011","100110011011","101010011100","101110101101","101110101100","100001111000","011001000101","010001000100","010000110011","010000110011","001100110011","010101000100","010101010101","010101000100","011101000100","011101000100","011101000100","011101000100","011000110100","011000110011","011000110011","011101000100","100001010101"),
		("101110111101","101110111101","101110111101","101010011011","100110011011","100110011011","101010101100","101110101101","101110101100","100001111001","010101000100","010101000100","010101000100","010000110011","010000110011","010101000100","010101010101","010101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","100001010101"),
		("101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010101100","101110101101","101110101101","100001111001","010100110100","010001000100","010101000100","010101000100","010000110100","010101000100","011001010101","011001010101","011101000100","011000110011","011000110010","011000110010","011000110011","011000110011","011000110011","011000110011","011101000101"),
		("101010101100","101110101101","101010011100","100110011011","100110011011","100110011011","101010101100","101010101100","101010101100","100001111000","010000110011","010000110011","010000110011","010000110011","010000110100","010101000101","011001010101","011001010101","011000110011","011000110010","010100100010","011000100010","011000110011","011000110011","011000110011","011000110011","011100110100"),
		("101010011100","101010101100","100110011011","100010001010","100110001010","100110001010","100110011011","101010011011","100110011011","011101100111","010000110011","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010101","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100110010"),
		("100110001010","100110001010","100001111001","100001111000","100001111001","100001111001","100010001010","100110001010","100110001010","011001010110","001100110011","001100100011","001100100011","001100110011","001100110011","010000110100","010101000100","010101000100","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010"))
	-- 11
	,

		(	("101010011100","101010101100","101010101100","101010101100","101010101100","101010011011","101010011011","100110011010","100110011011","100010001001","100001100111","100001010101","011000110011","010100100010","010100110010","011000110011","011000110011","011000110010","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011000110011","010100110010"),
		("101110101100","101110101101","101110101100","101110101101","101010101100","101010101100","101010101100","101010011011","101010011011","100110001001","100101100111","100001000101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000101","011101000101","011101000101","011101000101","011101000100","011000110011"),
		("101110101100","101110101100","101110101100","101110101100","101010101100","101010101100","101010011100","101010011011","101010011011","100101111001","100001010110","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001000101","100001000101","011101000101","011000110011"),
		("101110101101","101110101101","101110101101","101110101101","101110101101","101110101100","101010101100","101010101100","101010011011","100101111000","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001010110","011101000101","011000110011"),
		("101010101100","101010011100","101010011011","101010011100","101010011011","101010011011","100110001010","100110001010","100110001010","100101111000","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000100","100001000101","100001010110","100001000101","011000110100"),
		("100110001010","100110001011","100110011011","100110001011","100110001010","100110001010","100010001010","100001111001","100001111001","100001111001","100001010110","011100110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001000101","011100110100"),
		("100110001011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001","100101111000","100001010101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","011101000100"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100101111000","100001000101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001010110","100001010110","100001000101"),
		("100110011011","100110011011","100110011011","100110001010","101010011011","101010011011","100110011011","100110011011","100110001001","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","101010011011","101010011011","100110001010","100001111001","011101010101","011000100010","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001010","100110001010","101010011011","101010011011","100010001001","100001101000","011000110011","010100100010","011000110011","011000110011","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110010","011000110011","011101000100","011101000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100110001010","101010011011","100010001010","100001111001","011101010101","010100100010","010100110011","011000110011","011000110011","011000110011","010100110011","010000100010","010100100010","010100100010","010100110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110"),
		("100110001010","101010011011","101010011100","100110011011","100110001010","100001111001","100010001001","100110001010","100010001010","100010001001","100001100111","011000110100","011000110100","011000110011","011000110011","011000110100","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000101","100001010110","100001010110"),
		("101010011011","101010011011","101010011011","101010011100","100010001001","100001111001","100001111001","100010001001","100010001010","100010001001","100101100111","100001010101","011101000100","011000110011","011000110100","011000110100","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100001010110","100001010110"),
		("101010101100","101010101100","101010011100","101010011011","100010001001","100001111001","100001111001","100010001001","100010001010","100101111001","100101100111","100001010101","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101010101100","101110101100","101010101100","101010011011","100010001001","100001111001","100001111001","100010001001","100010001010","100101111000","100001010110","011000110100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","100010001001","100010001001","100010001010","100101110111","011101000100","011101000101","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001010101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011011","101010011011","100110001011","100110001010","100010001001","100010001001","100001010101","011100110100","100001000101","100001010110","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101010011100","101010011100","101010011011","101010011011","100110011011","100110011010","100110001001","100001111001","100001111001","011101010101","011000110100","011100110100","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","100001000101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111001","100001100111","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001000110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111001","100001111000","100001010101","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","011101000100","100001000101","100001000101","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101010101100","101010011100","100110001010","100001111001","100001111001","100001111001","100101100111","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","101110101100","100110001010","100001111001","100010001010","100110001010","100101100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110111101","101010101100","100110001010","100001111001","100010001001","100110011010","100101100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110101101","101010011100","100110001010","100010001001","100010001010","101010011011","100110001001","011101000100","011000110011","011000110011","011000110010","011000110010","011000110010","010100100010","010100100010","011000110011","011000110011","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010101100","100110001010","100110001010","100110001010","101010011011","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","011000110010","011000110011","011000110011","011000110100","011101000100","011101000100","100001000101","100001000101","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001001","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","100001000101","100001000101","100001000101","100001000101"),
		("101110111101","101110101101","101110101101","101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010001010","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011100110100","011101000100","011101000100","100001000101","100001000101"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010011100","100110001010","100110001010","100110011011","101010101100","101010101100","101010011011","100001100110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011000110100","011101000100","011101000100","011101000100","011101000101","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101110111101","101010011011","100110001010","100110001010","101010011011","101010101100","101010101100","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000101","011101000101","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100110001010","101010011011","101010011100","101010011100","101010101100","100101111000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101010101100","101010011011","100001100111","011000110100","011000110011","011000100010","011000110011","011000110011","011000110011","011000110100","011101000100","011100110100","011000110011","011000110011","011100110100","011101000100"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010101100","101110101101","101110101100","101010101100","101010101100","101110101100","101010011011","100101111000","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","101010011011","101010101100","101110101100","101010101100","101010101100","101010101100","101010101100","101110101100","101010101100","100001111000","011101000100","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110"),
		("101110111101","101110111110","101110111110","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","101110101101","101110101101","101110101100","101110101100","101110101101","101010101100","100001101000","011000110011","100001010101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011011","101110101101","101110101101","101110101101","101110101100","101010101100","101010011011","011101100110","011000110011","011000110011","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101"),
		("101110111101","101110101101","101110101101","101110101100","101010011011","100110011011","100110011011","101010011011","101110101100","101010011100","101010011010","100001111000","011101010110","011001000100","011000110011","011000110011","011101000100","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100"),
		("101110111101","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","101010011011","100110001010","011101100110","011001000100","011000110011","011000110011","011000110011","011000110011","011000110011","100001010110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100001111000","011001010110","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","100101100110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101110111101","101110101101","100110011011","100001111000","011001010101","010100110011","010100110011","010100110011","010100110011","010000100010","010000100010","010000100010","010100100010","010100100011","011001000100","100101100111","011101010110","010100110011","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101010011100","100001111000","011001010101","010100110011","010100100010","010000100010","010000100010","010101000100","010100110011","010000110011","010000110011","010101000100","010101000100","010101000100","011101100110","100101111000","011101100110","010100110011","010000100001","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("100110001001","011001010101","011000110011","010100110011","010000100010","010000100001","001100100001","001100100001","010000110011","010000110011","010000110011","010000110011","010000110100","010101000100","010101000101","011101100110","011101100111","011101100110","011001000100","010000100001","010000100010","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("011001000100","010100110011","010100100010","010000100010","001100100001","001000100001","001000010001","001000010001","010000100010","010101000101","010101000100","010000110011","010000110011","001100110011","010000110100","011001010110","010101000100","011101100110","011001010101","010000100010","010000100001","010100100010","010100110011","011000110011","011000110011","011000110011","011000110011"),
		("010100110011","010000100010","001100100001","001000100001","001000010001","001000010001","001000010001","001000010001","001100110010","010101000100","010000110100","010001000100","010000110100","010000110011","010000110011","011001010101","010101000101","011101100110","011101100110","010100110011","010000100001","010000100001","010100100010","011000110011","011000110011","011000110011","011000110011"),
		("010000100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100100010","010100110100","010000110011","010000110100","010000110100","010000110100","010001000100","011001010110","011001010101","011101100111","100001111001","011101100111","010100100010","010100100010","010100100010","011000110011","011000110011","011000110011","011000110011"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100110010","010100110100","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010110","011101100111","100001111000","100001111001","011001000100","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","010000110011","001100110011","001100110011","001100110011","010000110011","010000110100","011001010101","011001010101","011001010110","011101100110","100001111000","011101100111","010100110010","010100100010","010100100010","010100100010","010100100010","010100110010"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","001100110011","001100100010","001100100010","001100100010","001100100011","010000110011","010101000100","010101000100","011001010101","010101010101","011101100110","011101100111","010100110100","010100100010","010100100010","010100100010","010100100010","010100100010"))
	-- 12
	,

		(	("101010011100","101010101100","101010101100","101010101100","101010101100","101010011011","101010011011","100110011010","100110011011","100010001001","100001100111","100001010101","011000110011","010100100010","010100110010","011000110011","011000110011","011000110010","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011000110011","010100110010"),
		("101110101100","101110101101","101110101100","101110101101","101010101100","101010101100","101010101100","101010011011","101010011011","100110001001","100101100111","100001000101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000101","011101000101","011101000101","011101000101","011101000100","011000110011"),
		("101110101100","101110101100","101110101100","101110101100","101010101100","101010101100","101010011100","101010011011","101010011011","100101111001","100001010110","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001000101","100001000101","011101000101","011000110011"),
		("101110101101","101110101101","101110101101","101110101101","101110101101","101110101100","101010101100","101010101100","101010011011","100101111000","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001010110","011101000101","011000110011"),
		("101010101100","101010011100","101010011011","101010011100","101010011011","101010011011","100110001010","100110001010","100110001010","100101111000","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000100","100001000101","100001010110","100001000101","011000110100"),
		("100110001010","100110001011","100110011011","100110001011","100110001010","100110001010","100010001010","100001111001","100001111001","100001111001","100001010110","011100110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001000101","011100110100"),
		("100110001011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001","100101111000","100001010101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","011101000100"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100101111000","100001000101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001010110","100001010110","100001000101"),
		("100110011011","100110011011","100110011011","100110001010","101010011011","101010011011","100110011011","100110011011","100110001001","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","101010011011","101010011011","100110001010","100001111001","011101010101","011000100010","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001010","100110001010","101010011011","101010011011","100010001001","100001101000","011000110011","010100100010","011000110011","011000110011","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110010","011000110011","011101000100","011101000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100110001010","101010011011","100010001010","100001111001","011101010101","010100100010","010100110011","011000110011","011000110011","011000110011","010100110011","010000100010","010100100010","010100100010","010100110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110"),
		("100110001010","101010011011","101010011100","100110011011","100110001010","100001111001","100010001001","100110001010","100010001010","100010001001","100001100111","011000110100","011000110100","011000110011","011000110011","011000110100","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000101","100001010110","100001010110"),
		("101010011011","101010011011","101010011011","101010011100","100010001001","100001111001","100001111001","100010001001","100010001010","100010001001","100101100111","100001010101","011101000100","011000110011","011000110100","011000110100","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100001010110","100001010110"),
		("101010101100","101010101100","101010011100","101010011011","100010001001","100001111001","100001111001","100010001001","100010001010","100101111001","100101100111","100001010101","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101010101100","101110101100","101010101100","101010011011","100010001001","100001111001","100001111001","100010001001","100010001010","100101111000","100001010110","011000110100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","100010001001","100010001001","100010001010","100101110111","011101000100","011101000101","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001010101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011011","101010011011","100110001011","100110001010","100010001001","100010001001","100001010101","011100110100","100001000101","100001010110","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101010011100","101010011100","101010011011","101010011011","100110011011","100110011010","100110001001","100001111001","100001111001","011101010101","011000110100","011100110100","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","100001000101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111001","100001100111","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001000110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111001","100001111000","100001010101","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","011101000100","100001000101","100001000101","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101010101100","101010011100","100110001010","100001111001","100001111001","100001111001","100101100111","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","101110101100","100110001010","100001111001","100010001010","100110001010","100101100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110111101","101010101100","100110001010","100001111001","100010001001","100110011010","100101100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110101101","101010011100","100110001010","100010001001","100010001010","101010011011","100110001001","011101000100","011000110011","011000110011","011000110010","011000110010","011000110010","010100100010","010100100010","011000110011","011000110011","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010101100","100110001010","100110001010","100110001010","101010011011","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","011000110010","011000110011","011000110011","011000110100","011101000100","011101000100","100001000101","100001000101","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001001","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","100001000101","100001000101","100001000101","100001000101"),
		("101110111101","101110101101","101110101101","101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010001010","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011100110100","011101000100","011101000100","100001000101","100001000101"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010011100","100110001010","100110001010","100110011011","101010101100","101010101100","101010011011","100001100110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011000110100","011101000100","011101000100","011101000100","011101000101","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101110111101","101010011011","100110001010","100110001010","101010011011","101010101100","101010101100","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000101","011101000101","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100110001010","101010011011","101010011100","101010011100","101010101100","100101111000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101010101100","101010011011","100001100111","011000110100","011000110011","011000100010","011000110011","011000110011","011000110011","011000110100","011101000100","011100110100","011000110011","011000110011","011100110100","011101000100"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010101100","101110101101","101110101100","101010101100","101010101100","101110101100","101010011011","100101111000","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","101010011011","101010101100","101110101100","101010101100","101010101100","101010101100","101010101100","101110101100","101010101100","100001111000","011101000100","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110"),
		("101110111101","101110111110","101110111110","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","101110101101","101110101101","101110101100","101110101100","101110101101","101010101100","100001101000","011000110011","100001010101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011011","101110101101","101110101101","101110101101","101110101100","101010101100","101010011011","011101100110","011000110011","011000110011","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101"),
		("101110111101","101110101101","101110101101","101110101100","101010011011","100110011011","100110011011","101010011011","101110101100","101010011100","101010011010","100001111000","011101010110","011001000100","011000110011","011000110011","011101000100","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100"),
		("101110111101","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","101010011011","100110001010","011101100110","011001000100","011000110011","011000110011","011000110011","011000110011","011000110011","100001010110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100001111000","011001010110","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","100101100110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101110111101","101110101101","100110011011","100001111000","011001010101","010100110011","010100110011","010100110011","010100110011","010000100010","010000100010","010000100010","010100100010","010100100011","011001000100","100101100111","011101010110","010100110011","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101010011100","100001111000","011001010101","010100110011","010100100010","010000100010","010000100010","010101000100","010100110011","010000110011","010000110011","010101000100","010101000100","010101000100","011101100110","100101111000","011101100110","010100110011","010000100001","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("100110001001","011001010101","011000110011","010100110011","010000100010","010000100001","001100100001","001100100001","010000110011","010000110011","010000110011","010000110011","010000110100","010101000100","010101000101","011101100110","011101100111","011101100110","011001000100","010000100001","010000100010","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("011001000100","010100110011","010100100010","010000100010","001100100001","001000100001","001000010001","001000010001","010000100010","010101000101","010101000100","010000110011","010000110011","001100110011","010000110100","011001010110","010101000100","011101100110","011001010101","010000100010","010000100001","010100100010","010100110011","011000110011","011000110011","011000110011","011000110011"),
		("010100110011","010000100010","001100100001","001000100001","001000010001","001000010001","001000010001","001000010001","001100110010","010101000100","010000110100","010001000100","010000110100","010000110011","010000110011","011001010101","010101000101","011101100110","011101100110","010100110011","010000100001","010000100001","010100100010","011000110011","011000110011","011000110011","011000110011"),
		("010000100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100100010","010100110100","010000110011","010000110100","010000110100","010000110100","010001000100","011001010110","011001010101","011101100111","100001111001","011101100111","010100100010","010100100010","010100100010","011000110011","011000110011","011000110011","011000110011"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100110010","010100110100","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010110","011101100111","100001111000","100001111001","011001000100","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","010000110011","001100110011","001100110011","001100110011","010000110011","010000110100","011001010101","011001010101","011001010110","011101100110","100001111000","011101100111","010100110010","010100100010","010100100010","010100100010","010100100010","010100110010"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","001100110011","001100100010","001100100010","001100100010","001100100011","010000110011","010101000100","010101000100","011001010101","010101010101","011101100110","011101100111","010100110100","010100100010","010100100010","010100100010","010100100010","010100100010"))
	-- 13
	,

		(	("101010011100","101010101100","101010101100","101010101100","101010101100","101010011011","101010011011","100110011010","100110011011","100001111001","100001100111","011101000100","011000110011","010100110010","010100110011","011000110011","011000110011","011000110010","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011100110100","010100100010","010100100010"),
		("101110101100","101110101101","101110101100","101110101101","101010101100","101010101100","101010101100","101010011011","101010011011","100110001001","100101100111","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000101","011101000101","011101000101","011101000100","011000110011","011000110010"),
		("101110101100","101110101100","101110101100","101110101100","101010101100","101010101100","101010011100","101010011011","101010011011","100101111001","100001010110","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001000101","100001000101","100001000101","011000110011","010100100010"),
		("101110101101","101110101101","101110101101","101110101101","101110101101","101110101100","101010101100","101010101100","101010011011","100101111000","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001000101","100001000101","011101000101","011000110011","010100100010"),
		("101010101100","101010011100","101010011011","101010011100","101010011011","101010011011","100110001010","100110001010","100110001010","100101110111","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001000101","011000110011","011000110011"),
		("100110001010","100110001011","100110011011","100110001011","100110001010","100110001010","100010001010","100001111001","100001111001","100101100111","100001000101","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001010110","011000110011","011000110011"),
		("100110001011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001100110","011101000100","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100001000101","100001000101","100001010110","011100110100","011000110011"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001010110","011100110100","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","100001000101","100001000101","100001000101","100001010110","011101000101","011000110011"),
		("100110011011","100110011011","100110011011","100110001010","101010011011","101010011011","100110011011","100110011011","100101111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","100001000101","100001000101","100001000101","100001000101","100001010110","100001010110","011101000100"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","101010011011","101010011011","100110001010","011101010101","010100100010","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","011101000100","100001000101","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001010","100110001010","101010011011","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100110010","011000110011","010100110010","010100100010","011000110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100110001010","101010011011","100101111000","011000110011","010100100010","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000101","100001010110","100001010110","100001010110","100001010110"),
		("100110001010","101010011011","101010011100","100110011011","100110001010","100001111001","100010001001","100110001010","100110001001","011101000101","011001000100","011101000100","011000110011","011000110011","011000110100","011000110011","010000100010","010100100010","010000100010","010100100010","010100110010","011000110011","011101000100","100001010110","100001010110","100001010110","100001010110"),
		("101010011011","101010011011","101010011011","101010011100","100010001001","100001111001","100001111001","100010001001","100010001010","100101111000","100001010101","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101010101100","101010101100","101010011100","101010011011","100010001001","100001111001","100001111001","100010001001","100110001010","100001010110","011100110011","011000110011","011000110100","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110100","011100110100","011101000101","100001010110","100001010110","100001010110","100001010110"),
		("101010101100","101110101100","101010101100","101010011011","100010001001","100001111001","100001111001","100010001010","100001101000","011101000100","011101000100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","100010001010","100001111000","011101000101","011101000101","100001010110","100001000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001000101","100001010101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011011","101010011011","100110001011","100110001010","100001100111","011100110100","011101000101","100001000101","100001000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","100001000101","100001010110","100001010110"),
		("101010011100","101010011100","101010011011","101010011011","100110011011","100110011010","100110001010","100001111000","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","100001000101","100001000101","100001000101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","100001000101","100001000101","100001000110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","100110011011","100110001001","100001111001","100001100111","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001000101","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101010101100","101010011100","100110001010","100001111001","100101100111","100001010110","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","101110101100","100110001010","100010001001","100101111000","100001010101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110111101","101010101100","100110001010","100010001001","100001111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001000110","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110101101","101010011100","100110001010","100010001001","100001111001","011000110100","011000110011","010100100010","011000110011","011000110011","011000110010","011000110010","011000110010","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010101100","100110001010","100110001010","100010001001","100001010110","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110010","011000110011","011101000100","011101000100","011101000100","011101000100","011101000101","100001000101","100001000101","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101110111101","101010011011","100110001010","100110001010","100110001010","100110001001","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","100001000101","100001000101","100001000101","100001000101"),
		("101110111101","101110101101","101110101101","101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","101010011011","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001000101"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010011100","100110001010","100110001010","100110011011","101010101100","100101100111","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011000110100","011101000100","011000110100","011101000100","011101000100","011101000100","011101000101","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101110111101","101010011011","100110001010","100110001010","101010011011","101010101100","100101111000","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100110001010","101010011011","101010011100","100101100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000101","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010011100","101110101101","101010011010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001000110"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010101100","101110101101","101110101100","100110001010","011101010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011100110100","011101000100","011101000101","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","101010011011","101010101100","101110101100","101010101100","101010101100","101010011100","101010011010","100001100111","011101000100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001010110"),
		("101110111101","101110111101","101110111110","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","101110101101","101110101101","101110101100","101110101101","101010011011","011101010101","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110101101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011011","101110101101","101110101101","101110101101","101010101100","100101111001","011001000100","011101000100","100001010110","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","100001000101","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101010101100","100110011011","100110011011","100110011011","101010011100","101010101100","101010011011","100110001010","011101010110","011000110011","011000110011","100001010101","100001000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","100001000101","100001010110","100001010110","100001010110"),
		("101110101101","101110101100","101110101101","101110101100","100110001011","100110001010","100110001001","100001111000","011101100110","011001000100","011000110011","011000110011","011000110011","011001000100","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010101","100001010110"),
		("101110111101","101110101101","101110101101","101010011010","011101100111","011001000101","011000110100","010100110011","010100110011","010100100011","010100110011","010100110011","010100110011","100001010101","100001010101","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101"),
		("101010011011","100001111000","011101010110","011000110100","010100110011","010000100010","010000100010","010000100010","010000100010","010100110010","010000100010","010100110011","010100110011","100101100110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100"),
		("011001000100","011000110011","010100100010","010000100010","010000100010","001100100001","001100100001","001100100001","001100100001","011001000100","010000100010","010000110011","010100110100","011001000101","011001000101","011001000100","011101010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100"),
		("010100110011","010000100010","010000100001","001100100001","001000100001","001000010001","001100100001","001100100001","001100100001","010000110011","010000110011","010000110011","010001000100","010101000100","010101000100","010101010101","011101100111","011001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100"),
		("010000100010","001100100001","001000010001","001000010001","001000010001","001000100001","001000010001","001000010001","001000010001","010000110011","010101000100","010000110011","010000110011","001100110011","001100110011","010101000101","010101000101","010100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010100110100","010000110100","010000110100","010000110100","010000110011","010000110011","010101000100","010101000101","010100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","010000110011","010000110011","010000110100","010000110011","010101000100","011001010101","010101000100","011000110011","011000110011","011000110010","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","010000110011","010000110011","010000110011","010000110011","010101000101","011001010101","010101000100","010100100010","011000110011","011000110011","011000100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010000110011","010000110011","001100110011","001100110011","001100110011","010000110011","010101000100","011001010101","010101000100","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100110010"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010000110011","001100100010","001100100010","001100100010","001100100011","001100110011","010000110100","010101000100","010000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010"))
	-- 14
	,

		(	("101010011100","101010101100","100101111000","011101000100","010100100010","010000100001","010000100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100010001","001100010001"),
		("101110101100","101010101100","100001100111","011000110010","010100100010","010000100001","010000100001","001100100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("101110101100","101010011011","100001100111","011001000100","010100100010","010100100010","010000100001","010000100001","001100100001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("101110101101","101110101101","101010011011","100101111000","011000110011","010100100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("101010101100","101010011100","101010011011","100001111000","011101000100","010100110010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100010","001100100001","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001"),
		("100110001010","100110001010","100110001010","100001111000","011101000101","010100100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100010","010100100010","010100100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001"),
		("100110001011","100110011011","100110001010","100001111001","100001010110","011000110010","010000100001","001100100001","001100100001","010000100001","010000100010","010000100010","010100100010","011000110011","011000110011","011000110011","011100110011","011100110100","011000110011","010100110011","010100100010","010000100010","010000100001","010000100001","001100100001","001100100001","001100100001"),
		("100110011011","100110011011","100110011011","100110001010","100101111001","011101000101","010100100010","010000100010","010100100010","011000110011","011000110011","011000110011","011000110100","011000110011","011100110100","011101000100","011101000100","011101000100","011101000100","011000110011","011000110011","010100100010","010100100010","010000100010","010000100010","010000100010","010000100001"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100101100111","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","011101000101","011101000101","011101000101","011101000100","011100110100","011000110011","010100100010","010100100010","010000100010","010000100010","010000100001"),
		("100110011011","100110011011","100110001011","100110001010","100110001010","100101100110","011101000100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000101","100001000101","100001000101","100001000101","100001000101","011101000101","011000110011","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001"),
		("100110011011","100110011011","100110001010","100110001010","100101111000","100001010101","011101000100","011101000100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100001000101","100001000101","100001000101","100001010110","011101000101","011000110011","011000110011","010100100010","010000100010","010000100010","010000100010","010000100001"),
		("100110011011","100110011011","100110011011","100110001010","100101110111","100001010101","011101000100","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001010110","100001010110","100001000101","011000110011","011000110011","010100100010","010000100010","010000100010","010000100010","001100100001"),
		("100110001010","101010011011","101010011100","100110011011","100101110111","100001010101","011101000100","011100110011","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001010110","100001010110","100001000101","011100110100","011000110011","010100100010","010000100010","010000100010","010000100010","001100100001"),
		("101010011011","101010011011","101010011011","101010011011","100101111000","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110100","011000110011","011000110100","011000110100","100001000101","100001010110","100001010110","100001010110","011101000100","011000110011","010100110010","010000100010","010000100001","010000100010","010000100010"),
		("101010101100","101010101100","101010011100","101010011011","100101111000","011101000100","011100110011","011100110011","011000110011","011000110011","011000110011","011000110011","011000110100","011000110100","011000110100","011100110100","100001000101","100001010110","100001010110","100001010110","100001000101","011100110100","010100100010","010000100010","010100100010","010000100010","010000100010"),
		("101010101100","101110101100","101010101100","101010011011","100101100111","011101000100","011000110011","011100110011","011000110011","011000110100","011000110100","011000110011","011000110100","011000110100","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","011101000101","011000110011","010100100010","010100100010","010100100010","010100100010"),
		("101010011100","101010011100","101010101100","101010011011","100001100110","011100110011","011000110011","011000110011","011000110011","011000110011","010100110010","010100100010","010100110010","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001000101","011000110011","010100110011","010100110011","010100110011"),
		("101010101100","101010101100","101010101100","100110001010","011101000100","011000110011","011000110011","011000110011","011000110010","010100100010","010100100010","010100100010","010100100010","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","011101000101","011000110011","011000110011","011000110011"),
		("101010011100","101010011100","101010011100","100110001010","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100110010","011000110011","011000110011","011000110011","011101000101","100001000101","100001010110","100001010110","100001010110","100001010111","100001000101","011000110100","011000110011","011000110011"),
		("101010101100","101010101100","101010101100","101010011100","100001100111","011000110011","010100110010","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010100100010","011000110010","011000110011","011000110011","011000110100","100001000101","100001010110","100001010110","100001010110","100001010111","100001010110","011101000100","011000110011","011000110011"),
		("101010101100","101010101100","101010101100","101010011100","100110001001","011000110100","011000110100","011000110011","011000110011","011000110100","011000110011","010100100010","010000100010","010100100010","010100110011","011000110011","011000110011","011000110011","011101000100","100001010110","100001010110","100001010110","100001010111","100001010110","011101000100","011000110100","011000110100"),
		("101110101101","101110101101","101110101101","101110101101","101010011011","100101100111","100001000101","011000110011","011000110011","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","100001000101","100001010110","100001010110","100001010110","100001010111","100001010111","100001000101","011101000100","011101000100"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","100101111000","011100110011","011000110011","011000110011","011100110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","100101010111","100001010110","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101010011100","100001010101","011101000100","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","100101010111","100101010111","100101100111"),
		("101110111101","101110111101","101110111101","101110101101","100001100111","011101000100","100001010110","011101000101","011000110100","011000110011","011000110011","011000110010","011000110011","011000110011","011000110010","011000110011","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100101010111","100101010111","100101010111"),
		("101110111110","101110111110","101110111110","101010011011","011101000100","011101000101","100001000101","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100101010111","100101010111","100101010111"),
		("101110101101","101110101101","101110101101","101010011011","100001010110","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100101010111","100101010111","100001010110"),
		("101110111101","101110101101","101110101101","101110101101","100110001001","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001000101","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","100101010111","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101010001010","011101000101","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000101","011101000101","100001000101","100001010110","100001010110","100001010110","100101010111","100101010111","100001010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101010011011","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110","100101010111","100101010111","100001010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100101100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010111","100101010111","100101010111","100001010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101100","100001100111","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","100101010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101100","100001100111","011000110011","011000110011","011000110010","011000110010","011000100010","010100100010","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010111","100001010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110001001","011101000100","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000101","100001000101","100001000110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111110","101110111110","101010101100","100110001010","100001100111","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110101101","101110111101","101110111101","101010011100","100110011011","100101111001","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","100001000101","100001000101","100001000101","100001010110","100001000101","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101010101100","100110011011","100110011011","100110001010","100001100110","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001000101","100001000101","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("101110101101","101110101100","101110101101","101110101100","100110001010","100110001010","100110001010","100101111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000100","011101000100","011101000100","100001000101","011101000101","100001000101","100001000101","100001010110","100001010110","100001010110","100001010101"),
		("101110101101","101110101101","101110101101","101110101100","100110001010","100110001010","100110001010","100101111001","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001000101"),
		("101110101101","101110101100","101110101101","101010101100","100110001010","100110001010","100110001010","101010011011","011101010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010101","100001010110","100001010110","100001000101"),
		("101110111101","101110111101","101110111110","101010011100","100110001011","100110001010","100110011011","101010101100","100101111000","010100100010","010100110011","010100110100","010100110100","010101000100","010101000100","011101010110","011101000101","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101010011011","100110001011","100110001010","101010011011","101110101100","100001101000","010000100010","010000110011","010000110100","010001000100","010101000100","010101000101","011101100111","011001010101","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","100110011011","100110011011","100110001010","101010011011","101010101100","100101111001","011001000101","010000110100","010000110011","001100110011","001100110011","010101000100","011001010101","010100110100","011000110011","011000110011","011000110011","011101000100","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110111110","101110101101","100110011011","100110011011","100110001010","101010011011","101110101100","100001111001","010100110100","010000110100","010000110100","010000110011","010000110011","010000110100","011001010101","010101000100","011000110011","011000110011","011000110011","011101000100","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110111101","101010101100","100110001010","100110001010","100110001010","101010011011","101010011010","011101100111","010000110011","010000110100","010000110100","010101000100","010000110011","010101000100","011001010110","010101000101","011000110011","011000110011","011000110011","011100110100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","100110001010","100001111001","100001111001","011101100111","011101010110","011001000100","010101000100","010000110011","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010101","011000110011","011000110011","011000110010","011000110011","011101000100","011101000100","011101000101","100001000101","100001000101","100001010110"),
		("100110001010","100110001001","011101100110","011001000100","010100110011","010000100010","010000100001","001100100001","010000110011","010000110011","001100110011","001100110011","001100110011","010000110011","010101000100","011001010101","011001000101","010100110011","010100100010","010100100010","010100110010","011000110011","011000110011","011000110100","011101000100","011101000100","100001000101"),
		("011001000101","010100110011","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000110011","001100100011","001100100010","001100100010","001100100010","001100110011","010000110011","010101000100","010101000100","010100100010","010100100010","010100100010","010100100010","010100100010","010100110010","011000110011","011000110011","011000110100","011101000100"))
	-- 15
	,

		(	("101010011100","101010101100","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111000","100001111001","100110001010","100110001010","100110001001","100001111001","100001111000","100010001001","100010001001","100110001010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001"),
		("101110101100","101110101100","101010101100","101110101100","101010101100","101010101100","101010101100","101010011100","101010101100","100110001010","100001111001","100001111001","100110001010","101010011011","100110001011","100110001010","100110001010","100110001010","101010011010","100110011011","101010011011","101010011011","101010011011","101010011011","100110001010","100010001001","100010001010"),
		("101110101100","101010101100","101010101100","101010101100","101010101100","101010011100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111000","100001100111","100001100111","100001111000","100101111000","100101111001","100110001001","100110001010","100110011010","101010011011","101010011011","101010011011","101010011011","100110001010","100010001010","100010001010"),
		("101110101101","101110101101","101110101100","101110101101","101010101100","101010101100","101010011010","100110001001","100101100111","100001010101","011101000100","011000110011","011000110011","011000110010","011000110011","011000110011","011101000100","011101000100","100001010110","100101111000","100110001001","100110001001","100101111001","100110001001","100110001010","100010001001","100010001010"),
		("101010011100","101010011011","101010011011","101010011011","100110001001","100101100110","100001010100","011101000011","100001000011","011101000011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","011000110011","011100110011","011101000011","011101000100","011101000100","011101000100","011100110100","011101000101","100101111000","100001111001","100001111001"),
		("100110001010","100110001010","100110001010","100001100111","100001010100","100001000011","011101000011","100001000100","100001010100","100001000011","011000110011","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","011101000100","011101000101","100001010110","011101010101"),
		("100110001010","100101111000","100101100101","011101000011","011101000011","100001000100","011101000011","011101000011","011101000011","011000110010","010100100010","010000100010","010000100001","010000100001","010000100001","010000100001","010000100001","010000100010","010100100010","010100100010","010000100010","010000100001","010000100001","011000110011","011000110011","011000110011","011000110011"),
		("100101110111","100101100101","011101000011","010100100010","010100100010","010100100010","010000100001","010000100010","010000100001","010000100001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100001","001100100001","010000100001","010000100010","010000100001","001100100001","001100100001","010000100001","010100100010","011000110011","010100100010","010000100010"),
		("100001010100","011101000011","010100100010","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100001","010000100010","010000100010","010000100001","001100100001","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","010100100010","010100100010","010000100001"),
		("011100110011","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010000100001"),
		("011000110010","010100100010","010000100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100010","010000100010","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010000100010","010000100001"),
		("010100100010","010100100010","010000100001","010000100001","010000100001","001100100001","001100100001","010000100001","001100100001","001100100001","010000100001","010000100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100100001","001100100001","010000100001"),
		("011000110011","010100100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001"),
		("011101000101","011000110011","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("100001010110","011000110011","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("100101111000","011000110011","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100001","010000100010","010000100010","010000100001","010000100001","010000100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("100110001010","100001010110","010100100010","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100010","010100100010","010100100010","010100100010","010100100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101010101100","100110001001","011000110100","010000100010","010000100010","010100100010","010100110010","010100110010","010100110010","011000110011","011000110011","011000110100","011000110100","011000110100","011000110011","010100110011","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001","001100010001"),
		("101010011100","101010001010","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011000110100","011000110011","011000110011","010100100010","010100100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001","001100010001"),
		("101010101100","100110001001","100001010101","011101000100","011101000100","011100110100","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011101000100","011100110100","011000110011","010100100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101010011100","100101100111","100001000101","011101000100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011000110011","010100100010","010000100010","010000100010","010000100001","010000100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101100","100101100111","011101000100","011101000100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","100001000101","100001000101","011000110100","011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101100","100101100111","011101000100","011101000100","011000110100","011000110011","011000110011","011100110011","011000110011","011100110011","011000110011","011000110100","011101000100","100001000101","100001000101","011100110100","011000110011","010100100010","010000100010","010000100010","010000100010","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101100","100101100110","011101000100","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","011101000100","011000110011","010100110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001"),
		("101010101100","100001010110","011100110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","011101000100","011000110011","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001"),
		("101010101100","100001010101","011000110011","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","011101000101","011000110100","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001"),
		("101010001010","011101000100","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","011101000100","011000110011","010100100010","010000100010","010000100010","010100100010","010100100010","010000100010","010000100010","010000100001","010000100001"),
		("100001101000","011000110011","011000110011","011000110011","011000110011","011000110011","010100110011","010100100010","010100100011","011000110011","011000110011","011000110011","011101000101","100001000101","100001000101","100001000101","011101000101","100001000101","011100110100","010100110010","010100100010","010100100010","010100100011","010100100010","010100100010","010000100010","010000100010"),
		("101010011011","011001000100","011000110011","011000110011","010100100010","010100100010","010100100010","010000100010","010100100010","010100100010","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","011101000101","100001000101","100001000101","011100110100","010100110011","010100110011","010100110011","010100110011","010100110011","010100110011","010100100010"),
		("101110101101","100001101000","010100100010","011000110011","011000110011","010100110011","010100100010","010100100010","010100100010","010100100010","010100110010","011000110011","011000110011","011100110100","100001000101","100001000101","011101000101","100001000110","100001000101","011101000100","011000110011","010100110011","010100110011","010100110011","010100110011","010100110011","010100110011"),
		("101110111101","101110101100","011101000101","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010000100010","010100100010","010100100010","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001000101","011101000101","011000110011","011000110011","011000110011","010100110011","010100110011","010100110011","010100110011"),
		("101110111110","101110101101","100001100110","011000110100","011000110100","011000110100","011000110011","010100110010","010100100010","010100100010","010100100010","010100110010","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001000101","100001000101","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111110","101110101100","100001010101","011000110011","011000110100","011000110100","011000110011","011000110011","011000110010","011000110011","011000100010","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","011101000101","011000110100","011000110011","011101000100","011100110100","011000110011","011000110100"),
		("101110111110","100101111001","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001000101","100001000101","100001010110","100001010110","011100110100","011100110100"),
		("101110101100","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100101010111","100001010110","100001000101","011000110011"),
		("100001100111","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","100001010101","100001000110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","011000110011"),
		("011100110100","011101000100","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","011101010101","011101000100"),
		("100001010110","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001000101","011101000100","011100110100","011101000101"),
		("101110101100","100001010110","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001010110","100001010110","100001010110","100001010111","100001010110","100001010110","011101000100","011000110011","011000110011","011101000100"),
		("101110101101","100110001001","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011000110011","011000110011","011000110011","011100110100","011100110100","011101000100","011101000100","100001010110","100001010110","100001010110","100001010111","100001010110","100001010110","011000110011","011000110011","011000110011","011100110100"),
		("101110111110","101010101100","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","010000100010","010000110011","010100110100","010101000100","010101000100","011001000100","100001100111","100001100111","100001010110","100001010110","100001010111","100001010111","100001010110","011000110100","011101000100","011101000101","100001000101"),
		("101110111101","101110101101","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010000110011","001100110011","010000110100","010101000100","010101000100","010101010101","011101100111","011101010110","100001000110","100001010110","100001010111","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","100101101000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","010101000100","010000110011","010000110011","001100110011","001100100011","010101000100","011001010101","010101000100","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110111110","101010011011","011101000100","011000110011","011000110010","010100100010","011000110010","010100100010","011000110100","010100110100","010000110100","010001000100","010000110011","010000110011","010001000100","011001010101","011001000100","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110111101","101010101100","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011001000100","010000110011","010000110011","010000110100","010000110100","010000110011","010101000100","011001010101","011001010101","100001010110","100001010110","100001010110","100001010110","100001000101","100001010110","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","100110011011","100001101000","011000110011","011000110011","011000110011","011000110011","011000110011","011001000100","010000110011","010000110011","010000110011","010000110011","010000110100","010101000100","011001010101","011101010101","100001000101","100001000101","100001010110","100001010110","011101000101","011101000101","100001000101","100001000101","100001010110"),
		("101010011011","101010011011","100110001010","100001111000","011001000100","010100110011","010100110011","010100100010","010100100010","010100110100","010000110011","001100110011","001100110011","001100110011","010000110011","010101000100","011001010101","011001010101","011101000100","011101000100","011101000101","011101000101","011101000100","011000110100","011101000100","011101000100","100001000101"),
		("100110001010","100110001010","100001111000","100001111000","011001000100","010100100011","010100100010","010000100010","010000100010","010000110011","001100100010","001100100010","001100100010","001100100011","001100110011","010000110100","010101000100","010101000100","011000110100","011000110100","011101000100","011001000100","011000110100","011000110011","011000110100","011000110100","011101000100"))
	-- 16
	,

		(	("101010011100","101010101100","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001","100001111001","100110001010","100110001010","100110001010","100010001001","100001111001","100010001001","100110001001","100110001010","100110001010","100110001010","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101110101100","101010101100","101110101100","101010101100","101010101100","101010101100","101010011100","101010011100","100110001010","100001111001","100001111001","100110001010","101010011011","100110011011","100110001010","100110001010","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100010001010","100010001010"),
		("101110101100","101010101100","101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100110001010","101010011011","100110011011","100110011011","100110001010","100110001010","101010011011","101010011011","101010011100","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010"),
		("101110101101","101110101101","101110101100","101110101100","101010101100","101110101100","101010101100","101010101100","101010011100","100110001010","100010001010","100010001010","100110011011","101010011011","101010011011","101010011011","101010011011","101010011011","101010101100","101010101100","101110101100","101110101100","101110101100","101110101100","100110001010","100110001010","100110001010"),
		("101010011100","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100110001010","100010001010","100010001001","100001111001","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010"),
		("100110001010","100110001010","100110001011","100110011011","100110011011","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100010001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010"),
		("100110001011","100110011011","100110011011","100110011011","100110011011","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100010001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100010001010","100010001010","100010001001","100001111001","100001111001","100001111001","100010001001","100010001001","100010001001","100001111001","100001111001","100001111001","100010001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010"),
		("100110011011","100110011011","100110011011","100110011011","101010011011","101010011011","100110011011","100110011011","100101111001","100001111000","100001100111","100001100111","100001100111","100001100111","011101010110","011101010101","100001010110","100001100111","100101111001","100110001010","100110011010","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010"),
		("100110011011","100110011011","100110011011","100110001011","100110001011","100110011010","100110001001","100001100110","100001000100","011101000011","011100110011","011100110011","011100110011","011000110011","010100100010","010100100010","011000110010","011000110011","011101000100","011101000101","100001100111","100110001010","100110001010","100110001010","100010001001","100010001010","100110001010"),
		("100110011011","100110011011","100110001010","100110001001","100101111000","100101100110","100101010101","011100110011","011000110011","011000110010","010100110010","011000110011","011000110011","011000110010","010100100010","010100100010","010100100010","010100100010","011000110011","011000110011","011101000100","100001010110","100001100110","100001100111","100001100111","100001111000","100110001010"),
		("100110001011","100110001010","100101111001","100101100110","100101100101","100101100101","011101000011","010100100010","011000110011","011100110011","011101000011","011101000011","011101000011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","011000110010","010100110010","011000110011","011100110100","011100110100","011000110011","100001010101","100101111001"),
		("100110001010","100101111000","100101010101","100101010100","100101010100","011100110011","010100100010","001100100001","010000100001","010000100001","010000100001","010000100001","010100100010","010100100010","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010100100010","010100100010","010100100010","011000110011","011101000101","100001100110"),
		("100110001001","100101100101","011101000011","011000110011","011000110010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010000100010","010000100010","010100100010","010100100010","010000100010","011000110011","011101000100"),
		("100101111000","100001010101","011100110011","010100100010","010100100010","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100010","010000100010","001100100001","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100001","010000100010","011000110100"),
		("100001010101","011000110011","010100100010","010100100010","010100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100010","010000100010","010100100010","010100100011","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","001100100001","001100100001","001100100001","010100100010"),
		("100001100111","010100110011","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100001","010000100010","010000100010","010000100001","010000100010","010000100001","001100100001","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100010001","001100100001"),
		("101010011011","011101000101","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001"),
		("100110011010","100001010110","011000110010","010100100010","010000100010","010000100001","001100100001","001100100001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001"),
		("101010011011","100001010110","011000110011","010100100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101010011011","100101111000","011000110011","010100100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101101","101010011011","100001010110","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010000100010","010000100010","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101101","101110101100","100101111001","011000110100","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010100100010","010100110011","010100110011","010100100011","010100100010","010000100010","010000100010","010000100010","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101101","101010101100","100101111000","011101000100","011000110011","010100110011","010100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011100110100","011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001"),
		("101110101101","101010001010","100001010101","011101000100","011000110100","011000110011","011000110011","011000110011","011000110100","011000110011","011101000100","011101000101","011101000101","100001000101","100001000101","100001000101","100001010101","011101000100","011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100010001","001100010001"),
		("101110101101","100101111000","011101000100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","100001000101","100001000101","100001000101","100001010110","100001000101","011000110100","010100110011","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001"),
		("101010101100","100001100111","011100110100","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","100001000101","100001010110","100001000101","011100110100","010100110011","010100100010","010100100010","010000100010","010000100001","001100100001","001100100001","001100100001"),
		("101010101100","100001100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001000101","100001010110","100001000101","011000110100","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001"),
		("101010101100","100101100111","011101000100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001000101","100001000101","100001010110","100001000101","011000110011","010100110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001"),
		("101010011011","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001010110","100001000101","011000110100","010100110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100010001"),
		("100110001001","100001010101","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011000110011","011000110011","011000110100","011101000101","100001000101","100001010110","100001000101","011000110100","011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001"),
		("100001010101","011101000100","011000110011","011000110011","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110100","011000110100","011000110011","011100110100","100001000101","100001000101","100001010110","100001000101","011000110100","010100110011","010100100010","010000100010","010000100010","010000100001","010000100001","001100100001","001100100001"),
		("011001000100","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000101","100001000101","100001000101","100001010110","100001010110","011101000100","010100110011","010000100010","010000100010","010000100010","010000100010","010000100010","010000100001","010000100001"),
		("100101111000","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010000100010","010100100010","010100100010","011000110011","011100110100","011101000101","100001000101","100001000101","100001000101","100001010110","100001010110","100001000101","011000110011","010000100010","010000100010","010100100010","010100100010","010000100010","010000100010","010000100010"),
		("101010011011","011001000100","010100100010","011000110011","011000110011","011000110011","010100100010","010000100010","010000100010","010000100010","010100100010","011000110011","011000110100","011101000101","100001000101","100001000101","100001010110","100001010110","100001010110","011101000101","011000110011","010100100010","010100100011","010100110011","010100100010","010100100010","010100100010"),
		("101010011011","011101010101","010100100010","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","011000110011","010100110011","010100100010","010100100010","011000110011","011101000101","100001000101","100001000101","100001010110","100001010110","100001010110","011101000100","010100110011","010100110011","010100110011","010100110011","010100110011","010100110011"),
		("101010001010","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","010000100010","010000100010","010100100010","010100100010","010100100010","011000110011","011100110100","100001000101","100001000101","100001010110","100001010110","100001010110","011101000101","011000110011","010100110011","010100110011","010100110011","011001000100","010100110011"),
		("100101110111","100001010101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010000100010","010100100010","010100110011","011000110011","011000110011","011101000101","100001010110","100001010110","100001010110","100001010110","100001000101","011000110011","010100110011","010100110011","010100110011","010100110011","011000110011"),
		("100001010110","100001010101","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011100110100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","011000110100","010100110011","010100110011","010100110011","011000110011","011000110011"),
		("100101100110","011101000101","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","011101000100","011000110011","011000110100","011000110100","011000110011","011100110100"),
		("100001010101","011101000100","100001010110","100001010110","100001000101","011000110011","011000110011","011000110011","011101000100","010100110011","010000100010","010100110011","010101000100","011001000100","011001000100","011101010101","100001100111","100001010110","100001010110","100001010110","100001010111","100001010110","011101000101","100001010110","100001000101","011000110011","011100110100"),
		("011100110100","011101000101","100001010110","100001010110","100001010110","011100110100","011000110011","011000110011","011000110100","010000110011","010000110011","010000110011","010001000100","010101000100","010101000100","011001100110","011101100111","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100101010111","100001010110","011101000100","011000110011"),
		("011000110100","011000110100","011000110011","011100110100","100001000101","011000110100","011000110011","011000110011","011000110011","011001000100","010101000100","010000110011","010000110011","001100110011","010000110011","011001010110","010101000100","011101010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","011101000100","011000110011"),
		("011100110100","011000110100","010100110010","010100100010","011000110011","011000110011","010100100010","010100100010","011000110011","011000110100","010000110011","010000110100","010000110100","010000110011","010000110011","011001010101","010101000100","011101010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","011101000100","011100110100"),
		("011101000101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100110100","010000110011","010000110100","010000110100","010000110011","010000110011","011001010101","011001010101","011101010110","100001000110","100001010110","100001010110","100001010110","100001000101","100001000101","011101000100","011101000100","100001010110"),
		("100001010101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100110100","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010101","100001010110","100001000101","100001000101","100001010110","100001010110","011101000101","011000110100","011000110011","011101000100","100001010110"),
		("011101000101","011000110011","011000110011","011000110011","011000110011","010100110011","010100100011","010000100010","010100110011","010100110011","001100110011","001100110011","001100110011","010000110011","010000110011","011001010101","011001010101","011101010101","011101000101","011101000100","011101000101","011101000101","011000110100","010100100010","011000110011","011000110011","011101000101"),
		("011001000101","010100100010","010100100010","010100100010","010000100010","010000100010","010000100001","010000100001","010000100010","010000110011","001100100010","001100100010","001100100010","001100110011","010000110011","010101000100","010101000101","011001000100","011000110100","011000110100","011101000100","011101000100","010100110011","010100100010","011000110011","011000110100","011101000100"))
	-- 17
	,

		(	("101010011100","101010101100","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001","100001111001","100110001010","100110001010","100110001010","100010001001","100001111001","100010001001","100110001001","100110001010","100110001010","100110001010","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101110101100","101010101100","101110101100","101010101100","101010101100","101010101100","101010101100","101010101100","100110001010","100001111001","100001111001","100110001010","101010011011","100110001011","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100010001010","100010001010"),
		("101110101100","101010101100","101010101100","101010101100","101010101100","101010101100","101010011011","101010001010","100101111001","100101100110","100101100101","100001010110","100101110111","100101111000","100101111000","100110001001","100110001010","100110001010","101010011011","101010011011","101010011100","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010"),
		("101110101101","101110101101","101110101100","101110101101","101010011011","100110001001","100001010110","100001010101","011101000100","011100110011","011101000011","100001010100","100001000100","100001000011","100001010100","100101100101","100101100110","100101100111","100101111000","100110001001","101010011011","101010101100","101110101100","101110101100","100110001010","100110001010","100110001010"),
		("101010011100","101010011100","101010011011","101010001010","100101100110","011101000011","010100100010","011000110010","011000110011","011100110011","100001000011","100001000011","011000110011","011100110011","100001000011","011101000011","011101000011","100001000100","100001010101","100101100110","100101110111","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010"),
		("100110001010","100110001010","100101111000","100101100101","100001010100","011000110010","010100100010","100001000100","100001000011","100001000011","100001000011","011000110011","011000110011","011000110011","010100100010","010000100001","010000100001","011000110011","011000110011","011101000100","100001010101","100101100110","100101111000","100010001001","100110001010","100110001010","100110001010"),
		("100110001011","100101111001","100101010101","100101010100","100001000100","011000110010","100001000100","100101010100","011100110011","011000110010","011000110010","010100100010","010000100010","010000100001","010000100001","001100100001","001100100001","010000100010","010100100010","010100100010","011101000100","100001010110","100101100111","100001100111","100001100111","100110001001","100110001010"),
		("100110001010","100101100110","100001000011","100001000100","011101000011","011101000011","100001000011","011101000011","010100100010","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010100110011","011000110011","011000110011","011000110100","011101000100","011101010110","100001111000"),
		("100101100110","011101000011","011000110011","010100100010","010100110010","010100100010","010000100010","010000100001","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100001","010100100010","011000110011","011101000100","011000110011","010100110010","100001010101"),
		("100101100101","011000110010","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100100010","011000110011","011101000101","011101000101","010100110011","010100110011","011101000101"),
		("100001010100","011000110010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","010000100010","010000100010","010000100010","010100110011","011000110011","011101000100","011101000100","011101000100","011000110011","011000110011","011101000101"),
		("011000110011","010100110010","010000100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","010000100010","010100100010","010100100010","010100100010","010000100010","010000100010","010100100010","010100110010","010100100010","010100100010","011000110011","011000110011","011000110100","011000110011"),
		("011000110010","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100110011","011000110011","011000110011","011000110011"),
		("010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100100010","010100110011","010100110011","010100110011"),
		("010100100010","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100100010","010000100010","010000100010","010100100010"),
		("011000110011","010100100010","010100100010","010000100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100100010","010000100010","010000100001","010000100010"),
		("011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010100100010","010100100010","010100100010","010000100010","010000100010"),
		("011000110011","010100100010","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","001100100001","010000100001","010000100010","010100100010","010100110011","011000110011","011000110011","011000110011","010100110011","010000100010","010000100010"),
		("010100100010","010100100010","010100100010","010100100010","010100110011","010100110011","010100110011","010100110011","010100110011","010100110010","010100100010","010000100010","010000100010","010000100010","010100100010","010100110011","011000110011","011101000100","011101000101","011101000101","100001010110","100001010110","100001010110","100001010101","011000110100","010100100010","010000100010"),
		("010100100010","010100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001010110","100001010110","100101100111","100101100111","100101100111","100101100111","100101100111","100101100111","011101000101","010100110011","010100100010"),
		("010100100010","010100110011","011000110011","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011101000100","011101000101","100001010110","100001010110","100001010110","100001010111","100101100111","100101101000","100101101000","100101100111","100101100111","100101100111","100001010110","011000110011","010100110011"),
		("010100100010","011000110011","011000110011","011000110011","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011101000100","011101000100","011101000101","100001010101","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101100111","100101100111","100101100111","100001010110","011000110100","010100110011"),
		("010100100010","011000110011","011000110100","011000110100","011000110011","011000110100","011000110100","011000110011","011000110100","011000110100","011101000100","011101000100","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101100111","100101100111","100001010110","011000110100","010100110011"),
		("010100110011","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000101","100001000101","100001010101","100001010110","100101010111","100101010111","100101100111","100101100111","100101010111","100001010110","011000110100","011000110011"),
		("010100110011","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110100","011000110011","011101000100","011101000100","011101000101","100001000101","100001000101","100001000101","100001000101","100001000101","100001010110","100101010111","100101010111","100101010111","100101100111","100101010111","100001010110","011101000100","011000110011"),
		("011000110011","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","100001000101","100001000101","100001000101","100001010110","100001010110","100001010111","100101010111","100101010111","100101010111","100101010111","100101010111","100001010110","011000110100","011000110011"),
		("011000110011","011000110011","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","011101000100","011101000101","100001000101","100001010110","100001010110","100101010111","100101010111","100101010111","100101010111","100101010111","100101010111","100001010110","011000110100","011000110011"),
		("011000110100","011000110100","011000110100","011000110011","010100110011","010100110011","010100110011","010100110011","010100110011","011000110011","011000110100","011101000100","011101000101","011101000100","011101000100","100001000101","100001010110","100001010110","100101010111","100101010111","100101010111","100101010111","100101010111","100101010111","100001010110","011000110100","011000110011"),
		("011101000100","011101000100","011000110011","010100110011","010100100010","010100100010","010000100010","010000100010","010000100010","010100100010","010100110011","011000110011","011000110100","011000110011","011000110011","011100110100","011101000101","100001000101","100001010110","100001010110","100101010110","100101010111","100101010111","100101010111","100101010111","011101000100","011000110011"),
		("011101000101","011101000100","011000110100","011000110011","011000110011","011000110011","010100110011","011000110011","010100100010","010100100010","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001010110","100001010110","100101010111","100101010111","011101000100","011000110100"),
		("100001010101","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","011000110011","011000110011","011101000100","011000110011","011000100011","011000110010","010100110010","011000110011","011000110011","011000110100","011101000100","100001010110","100101010111","100101100111","011101000100","011101000100"),
		("100101100101","011101000100","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011000110011","100001000101","100001010110","011101000101","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001000101","100001010110","100101100111","100101101000","011101000101","100001010110"),
		("100001010101","011101000100","011000110011","011000110011","011000110011","010100100010","010100110010","010100100010","011000110011","011000110011","011000110011","011000110011","100001010110","100101010111","100101010110","011101000101","011000110011","011000110011","011000110100","011101000101","100001010110","100001010110","100101010111","100101101000","100101111000","100001010101","100101100111"),
		("100001010101","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","100001010110","100101100111","100101100111","100001010110","011101000101","011101000100","011101000101","100001010101","100101010111","100101100111","100101100111","100101111000","100101111000","100001010101","100001000101"),
		("011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110","100101100111","100101100111","100101100111","100001010110","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101111000","100101111000","100001010110","011101000101"),
		("011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100101100111","100101100111","100101100111","100101100111","100001010110","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101111000","100101111000","100001010111","100001010110"),
		("100001000101","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100101010111","100101100111","100101100111","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101100111","100001100111","100101111000"),
		("100001010110","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","100001000101","100101100111","100101100111","100101010111","100001010110","100001000110","100001010110","100001010110","100001010110","100001010110","100101010111","100101100111","100101100111","100101100111","100101111000","100110001010"),
		("100101111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110","100001010110","100001010110","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001010111","100101100111","100101100111","100101100111","100110001001","101010011011"),
		("100101111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011000110100","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100101100111","100101111001","100110001010","100110001010","101010011011"),
		("100110001001","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011000110011","010000100010","010100110011","010100110100","010101000100","010101000100","011001010101","100101111000","100001010110","100001010110","100001010110","100001010110","100001010111","100101111000","100110001010","101010011011","101010011011","101010101100"),
		("101010001010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100110011","010000110011","010000110011","010000110100","010001000100","010101000100","011001010110","011101100111","100001010110","100001000110","100001010110","100001010110","100101010111","100101111000","100110011011","101010101100","101010011100","101010101100"),
		("101010011010","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011001000100","010101000100","010000110011","010000110011","001100110011","001100100011","011001010101","010101000101","011101010110","100001010110","100001010110","100001010110","100101100111","100101111000","101010011011","101010101100","101010101100","101110101101"),
		("101010011011","100001010110","011000110011","011000110011","011000110011","011000110010","010100100010","010100100010","011000110011","011001000100","010000110011","010001000100","010000110100","010000110011","010000110011","010101010101","010101000101","011101010110","100001010110","100001010110","100001010110","100101100111","100110001001","101010011011","101010011100","101010101100","101110101100"),
		("100110001001","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","010000110011","010000110100","010000110011","010000110100","010000110011","011001010101","011001010101","100001010110","100001000110","100001010110","100001010110","100101101000","100001111001","101010011011","101010011100","101010011100","101110101100"),
		("011101010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010101000100","010000110011","010000110011","010000110011","010000110011","010000110100","011001010101","011001010101","100001010110","100001000101","100001000101","100001010110","100001111000","100001111001","101010011011","101010011011","101010011011","101110101100"),
		("011101000101","011101000100","011000110011","011000110011","011000110011","010100110011","010100100011","010100100010","010100110010","010100110100","001100110011","001100110011","001100110011","010000110011","010000110011","010101010101","011001010101","011101010110","011101000101","100001000101","100001010110","100001100111","100001111001","100110001010","100110001011","100110011011","101010011011"),
		("011000110100","010100110011","010100100010","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000110011","001100100010","001100100010","001100100010","001100100011","010000110011","010101000100","010101000100","011001010101","011101000100","011101010101","011101010101","011101010110","100001100111","100001111001","100001111001","100001111001","100010001001"))
	-- 18
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010011011","101010011100","101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001010","100110011011","101010101100","101010101100","101010101100","101010101100","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110011010","100110001010","100101110111","100101110111","100101111000","100101111000","100110001001","101010011010","100110001010","100110001010","100110001010","100110001010","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001010","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011011","100101100111","100001000011","011100110011","011000110010","011000100010","011000110010","011101000101","100101111000","101010011011","101010101100","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010001010","100001000100","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","100001010101","101010011011","101010101100","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","101010001010","100101100110","011100110011","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011000110011","100110001001","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","101010011011","101010001001","100001010100","011000110011","011101000100","011101000101","100001010101","100001010110","100101100110","100001010110","011000110011","100101111000","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100110001010","101010011100","101010011010","011101000011","011101000100","100001010101","100001010101","100101100110","100101100110","100101100110","100101100110","011101000100","100001100111","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100110001010","100110001010","101010001010","011101000100","011101000100","011101000101","011101000100","100001010101","100101100110","100101010110","100101100110","011101000101","100001111000","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","100010001001","100110001010","011101010101","011101000100","011101000100","011101000100","011101000100","100001010101","011101000101","100001010101","100001010110","100001111000","100110011011","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011010","101010011011","100001111001","100001111000","100001010110","011101000100","011101000100","011101000100","011101000100","100001010110","100101010110","100101010110","100101100110","100001111000","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100010001010","100110001010","100101111001","100001000101","011101000101","011101000101","011101000100","011101000100","100001010101","100101100110","100101100110","100101100110","100110001001","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","100001100110","011101000101","011101000100","011101000100","011101000100","100001010101","100101100110","100101100110","100101100111","100110001001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011100","101010011011","100110001010","100110001010","101010011011","101010011011","100110011011","100001111001","100001100111","011101000101","011101000100","011101000100","100001010101","100101010110","100101100110","100001111000","100001111001","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011011","100110011011","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100110001010","100001010101","011101000100","011101000101","100001010110","100101100110","100101100110","100001111000","100110001010","100110001010","100001111001","100110001010","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100110001010","101010011010","100001100110","100001010110","011101000101","100001010101","100001010110","100001010110","100001100111","011101100111","101010011010","100110001001","100001111001","100110001010","100001111001","100001111000","100001111000"),
		("100010001001","100110001010","101010011100","101010011100","100110011011","100110001010","100110001010","100010001001","100001111001","100001111001","100110001010","100110001010","011101010101","011001010101","011101000101","011101000101","100001010110","100001010110","100001100111","010000110011","010101000100","011101100110","100001100111","100001111000","100001111001","100001111001","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110011011","100110001010","100110001010","100110001001","100001111001","100110001001","101010011010","100110001001","011001010101","011001010101","011101010101","100001000101","100001010110","100001100111","011101100111","001100100010","001100100010","001100100010","010000100010","010101000100","011001010101","011101100111","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110011011","100110001010","100010001010","100110001010","100001111001","100001111001","100110001010","100101111000","011001010101","011001010101","011101010101","100001000101","100001010101","100001100111","011101100110","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","010000110011"),
		("101010011011","100110001010","100110001010","101010011011","100110011010","100010001001","100010001001","100110001010","100010001001","100001111000","011101100111","011101010101","011001010101","011001010101","011101000101","011101000100","011101000101","100101111001","011101100111","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010"),
		("101010101100","100110001010","100110001010","101010011011","100110001010","100010001001","100001111001","100010001001","100101111001","011101010101","010000100010","010100110011","011101010110","011001010101","011101000101","011101000100","100001100111","100001111001","010000110100","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110011010","100110001010","100110011010","100110001010","100110001010","100001111001","100010001001","100001111000","011001000100","010000100010","001100100001","010000110011","100001100111","011101100111","100001010110","100001010110","100001111000","011001010110","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001010","100110001010","100110001001","100010001001","100001111000","100001100110","011000110100","001100100001","001100100001","001000100001","001100100010","100001100111","011101100111","011001010101","011001010101","011001000101","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","101010011011","100110001010","100001111001","100001111001","011101010110","010000100010","001100100010","001000100010","001000100010","001000100010","001000100001","011101010110","011101100111","010101000101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","101010011011","101010011011","100110001001","100101111001","010101000100","001100100001","001000100010","001000100010","001000100001","001000100001","001000100001","010101000101","011001010110","010101000100","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("101010011100","101010011011","101010011011","100110011010","100101111001","010101000100","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010"),
		("101010011011","101010011011","101010011011","101010011010","100001111001","011001000101","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010000110100","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010"),
		("101010101100","101010101100","101010011011","100110001001","100001111001","011101010110","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010000110011","010101000100","010000110100","001100100010","001100100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","101010011100","100110001001","100001111000","100001111001","011101100111","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010000110011","010001000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100010","001000100010"),
		("100110001010","100110001010","100110001001","100110001001","100001111001","011101100111","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","001100110011","010000110100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010"),
		("100110001010","100110001001","101010011010","101010011010","100001111001","011101100111","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","001100110011","010000110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010"),
		("100110001010","100110001010","101010011011","100110011010","100001111001","100001111000","010000110011","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","001100110011","010000110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100010"),
		("100110001010","100110001010","100110011010","100110011010","100001111001","100001111000","011001010101","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","001100100010","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001001","100110001010","100010001001","100001111000","011101100110","001100100010","001000100001","001000100001","001000100001","001000010001","001100110011","001100100010","001100110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000010001","001000100001","001000100010"),
		("101010011011","101010011011","100110001001","100010001001","100010001001","100001111000","011001000100","001000100001","001000010001","001000010001","001000010001","001000010001","001100110011","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","000100010001","001100110010","001000100010"),
		("101010011100","101010011011","100110001010","100110001001","100001111001","100001111000","010000110011","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000010001","001000010001","001000100001","001000100001"),
		("100110001010","100110001010","100110001010","100001111000","100101111000","011101010110","010000100010","001000100001","001000010001","001000010001","001000010001","001000010001","001100110010","001100100010","001100100010","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","000100010001","001000010001","001000010001","001000100001"),
		("100110001010","100110001010","100101111000","100001010110","100001010110","100001010101","010000110011","001100100001","001000010001","001000010001","001000100001","001000100001","001100110010","001100100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000010001","000100010000","001000010001","001000100001","001000100001"),
		("100110001010","100110001001","011101010101","100001000101","100001010110","100001010110","010100110011","001000100001","001000010001","000100010001","001000100001","001000010001","001100110011","001100100010","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100001","001000010001","000100010000","000100010000","001000010001","001000100001","001000100010"),
		("100110011010","100101111001","011101000100","011101000100","100001010101","100001010110","011001000100","001000010001","000100010001","000100010001","001000100001","001000010001","001100110011","010000110011","010000110011","001100100010","001000100001","001000100010","001000100001","010000100011","010000100010","001100100001","001000010001","000100010001","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100001010110","011000110100","011101000101","100001010110","011101000100","001000010001","000100010000","000100010001","001000010001","001000010001","001100110011","010101000100","010101000100","010000110011","001000100001","001000100001","001000100001","010100110011","011100110100","011000110011","010100110011","001000100010","001000100001","001000100010","001000100010"),
		("100110001010","100110001001","100001111000","011101010110","011101000100","011101000100","010000100010","001000010001","001100110011","001000100010","000100010001","001000010001","001100110011","010101000100","010101000100","010000110100","001000100010","001000100001","001000010001","011000110011","011101000100","011101000100","011101000100","010000100011","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100001111001","100001111000","010000110011","001100010001","010000110011","011101100110","011101100111","001000100010","000100010001","001000010001","001100110011","010101000100","010101000100","010101000100","001000100010","001000010001","000100010000","010100110010","011101000101","011101010101","011101000101","010100110100","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","010101000101","001100110011","011101111000","100110001001","011101010110","001100100010","000100010001","000100010001","001100110011","010101000100","010101000100","010101000100","001000100010","000100010001","000100010000","001100100010","011101000100","011101000101","011101000101","011001000100","001000100010","001100100010","001100100010"),
		("011101100111","011101100111","100001100111","100001110111","100001100111","011101100111","100001111000","011101100110","010000110011","001100100010","000100010001","000100010000","001100110010","010100110100","010101000100","010101000100","001100100010","000100010001","000100010000","001000100001","010100110011","011101000100","011101000100","010100110100","001000100010","001000100010","001000100010"),
		("011101100110","011101100110","011101100110","011101100110","011101100110","011101100111","011101100111","010101000100","001100100010","001000100001","000100010001","000100010000","001100100010","010000110011","010000110100","010000110100","001100100010","000100010001","000100010000","000100010000","001100100010","010100110011","010100110011","010000100010","001000100001","001000100001","001000100010"))
	-- 19
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100010001001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","100110001001","100101100110","100101100110","100001100110","100001100110","100001111000","100110001010","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100010001001","100110001010","100110001001","011101000011","011000110010","010100100010","010100100010","010100100010","011000110011","100001100111","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100101111000","100101010101","011000110010","010000100001","010000100001","010000100001","010100100010","010100100010","011000110011","100101111000","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110011011","100110001001","100101010101","011101000011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000100010","011101010110","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001010","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011100","101010011010","100001010100","011000110010","011101000100","011101000101","100001010101","100001010101","100001010110","100001010110","011000110100","011101010110","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011010","011101000100","011000110011","100001010101","100001010101","100001010110","100101100110","100101100110","100101100110","100001000101","011101010110","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011100","101010011010","011101000100","011100110100","011101000101","011101000100","100001010101","100101100110","100101100110","100101100110","100001010101","011101010110","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010101100","101010011011","011101010101","011101000100","011101000100","011101000100","011101000100","100001010101","011101000101","011101000101","100001010101","100110001001","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100110001010","101010011011","101010011011","101010101100","100110001001","100001010101","011101000101","011101000101","100001010101","011101000100","100001010101","100101010110","100001010110","100001100110","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010101100","100101111000","100001000100","100001000101","011101000101","011101000101","011101000100","100001010101","100101100110","100101100111","100101100111","101010011010","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","100010001001","100110001010","101010011011","100110001001","100001010110","011101000101","011101000100","011101000100","011101000100","100001010101","100101100110","100101100110","100101111000","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011010","101010011011","100001111001","100001111001","100010001001","100001111001","100110001001","100001100111","011101000100","011101000100","011101000100","100001010110","100101010110","100101100111","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100010001010","100110001010","101010011010","100110001010","100010001001","100110001010","100001100111","011101000100","011101000101","100001010101","100101100110","100101100110","100001111000","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011011","100010001001","100110001001","100001010110","011101000100","011101000100","011101000100","100001010110","100101010110","100001101000","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011100","101010011011","100110001010","100110001010","101010011011","101010011011","100110011011","100010001001","100001111000","100001111000","100001010110","011101000100","011101000100","011101000100","100001010110","100001010110","011101010110","011001010110","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011011","100110011011","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100110001010","100101111000","100001010101","011101000101","011101000100","100001010101","100101100110","100101010111","011101010110","001100100011","010101000100","100001111000","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100001111000","100001100111","100101100111","100001010110","011101010101","011101000100","100001010101","100001010110","100001100111","011001010101","001100100010","001100100010","001100100010","010100110100","011101010110","100001111000","100001111001"),
		("100010001001","100110001010","101010011100","101010011100","100110011011","100110001010","100110001010","100010001001","100001111000","011101010110","010100110011","010100110011","011101010110","011001010101","011101010101","011101000101","011101000100","011101010101","100101111000","010101000100","001100100010","001100100010","001000100010","001000100001","001000100001","001100100010","010101000100"),
		("100010001010","100001111001","100110011011","101010011011","100110011011","100110001010","100101111001","011101010110","010100110011","010000100010","001100100001","010000110011","011001010101","011001010101","011101010101","011101000100","011101010101","100001111000","100110001001","010000110100","001100100010","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001"),
		("100110011011","100010001001","100110001010","101010011011","100110001010","011101100111","011001000100","010000100010","001100100010","001000100010","001000100001","001100100010","011001010101","011001010101","011101100110","100001010110","100101111000","100110001001","011001010101","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100110001010","101010011011","100110001001","010000110011","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","011001010101","011001010101","011001010110","011001010101","011001010110","011001010110","001100110011","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010"),
		("101010101100","100110001010","100110001010","101010011011","100001111001","010000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","011001010101","011001010101","010101000101","010101000101","010101000100","001100100010","011001000100","011001000100","010100110011","001100100010","001000100010","001000100010","001000100010","001000100010"),
		("100110011010","100110001010","100110011010","100110001010","100001111000","001100100010","001000100010","001000100010","001000100001","001000100001","001100100001","001100100001","010000110011","011101100110","010101000101","011001000101","010101000101","010000110011","010000110011","100001010101","100001000101","011101000101","011001000100","001100100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001010","100110001010","100110001001","100001111000","001100100010","001000100010","001000100001","001100100001","001100100001","001000100001","001000100001","010000110011","100001100111","011001010101","010101000100","010101000100","001100110011","010101000100","100001010101","011101000101","011101010101","011101000100","001100100010","001000100010","001000100010","001000100010"),
		("100110001010","101010011011","100110001010","100010001001","011101100111","001100100010","001000100001","001100100010","001000100010","001000100010","001000100010","001000100001","010101000100","100001111000","011001010101","010101000100","010000110011","001100100010","011001000100","100001000101","100001000101","100001010101","011101000100","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","101010011011","101010011011","100110001001","011101100111","001100100010","001100100001","001000100010","001000100010","001000100001","001000100001","001000100001","010000110011","011101100110","010101000101","010001000100","010000110011","001100100010","010000100010","011100110100","011101000101","100001010101","011101000100","001100100010","001000100010","001000100010","001000100010"),
		("101010011100","101010011011","101010011011","100110011010","011101100111","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010101000100","010001000100","010000110011","001000100010","001000100010","010100110011","011101000100","100001010101","011101000100","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","101010011011","101010011011","101010011011","011101100111","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010001000100","010000110100","001100110011","001000100010","001000100010","001100100010","011000110011","011101000101","011101000100","001100100010","001000100001","001000100010","001000100010"),
		("101010101100","101010101100","101010011011","100110001001","100001111000","001100100010","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110100","010000110100","001100100010","001100100010","001100100010","001000100010","001100100010","010100110011","010100110011","001100100010","001000100001","001000100010","001000100010"),
		("101010011011","101010011100","100110001001","100001111000","100001111000","010000100010","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010001000100","010000110011","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","001000100010","010000110011","001000100010","001000100010"),
		("100110001010","100110001010","100110001001","100110001001","100001111000","010000110011","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110011","010000110011","001100100010","001000100010","001000100010","001000100010","001000010001","001000100001","001000100001","001000100010","011001010101","001100100010","001000100001"),
		("100110001010","100110001001","101010011010","101010011010","011101100111","001100100010","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110011","001100110011","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000010001","001000010001","001000100010","001000100010","001000100010"),
		("100110001010","100110001010","101010011011","101010011010","011101010110","010000100010","011001000100","010000100010","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110011","001100100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110011010","100110011010","011101010110","100001010101","100001010101","011000110011","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110011","001100110010","001000100010","001000100001","001000010001","001000010001","000100010001","001000010001","000100010000","000100010000","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001001","100110001010","100001111000","100001010101","100001010101","011101000100","001100100010","001000100001","001000100001","001000010001","001100100010","010000110100","010000110011","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","001000010001","001000100001","001000100010"),
		("101010011011","101010011011","100110001001","100010001001","100001010110","011100110100","100001010101","100001000101","010000100010","001000010001","001000010001","001000010001","001100100010","010000110011","001100100010","001100100010","001000100001","001000010001","001000010001","000100010001","000100010000","001000100001","001100100010","001000010001","000100010001","001100110011","001000100001"),
		("101010011100","101010011011","100110001010","100110001001","100001100111","011101000100","011101000101","100001010101","010000100010","000100010001","001000010001","001000010001","001100110011","010000110011","001100100010","001100100010","001000100001","001000100001","000100010001","000100010000","000100010000","001000100001","001100110011","001000010001","001000010001","001000100001","001000100001"),
		("100110001010","100110001010","100110001010","100110001001","100001100111","011000110100","011101000100","011101000100","010000100010","001000100001","001000010001","001000010001","001100110010","010000110011","001000100010","001000100001","001000100001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001"),
		("100110001010","100110001010","100110001010","100110001001","100001111000","011001000100","010000100010","010000110010","011101100111","010000110011","001000010001","001000010001","001100110010","010000110100","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001010","100110001001","100110001001","011101100111","010000110011","011101100110","100101111000","001100110011","001000100001","001000100001","010000110011","010101000100","010101000100","001100100010","001000100001","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","000100010000","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001010","100110001001","100001111001","100001111001","100001111001","100110001001","100001110111","001100100010","001000100010","001000100010","010101000100","010101000101","010101000100","001100100010","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001001","100110001001","100001111000","100001111000","100001111000","100110001001","011101010110","001100110011","001100110011","001100100010","010101000100","010101000101","010101000100","001100110011","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100001111001","100001111000","100001111000","100001111000","100110001001","011001010101","001100100010","010000110011","001100110011","011001010101","010101000101","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100001111001","100001111000","100001111000","100001111000","100001111000","100101111001","010101000101","001100100010","001100100011","010000110011","010101010101","010101000101","010101000100","010000110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","100001110111","100001111000","100001111000","100001111001","010000110100","001000100010","001100100010","010000110100","010101000101","010101000101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001000100010"),
		("011101100111","011101100111","100001100111","100001110111","100001110111","100001111000","100001111000","011101100111","001100110011","001000100010","010000110011","010101000100","010101000100","010101000100","010101000101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("011101100110","011101100110","011101100110","011101100110","011101100110","011101100111","011101100111","011001010110","001100100010","001000100010","010000110011","010000110100","010000110100","010001000100","010101000100","010000110100","010000110011","001100100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010"))
	-- 20
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100001111001","100001111001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011010","101010001010","101010001010","101010011010","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010001010","100101100110","100001010100","100001000100","011101000100","011101010101","100001100111","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001001","100101100110","011000110010","010100100010","010100100010","010100100010","010100100010","011000110011","100001100111","100110001001","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110011010","100110001010","100101100110","100001000100","010100100010","010000100001","010000100001","010000100001","010000100001","010100100010","011000110011","100001111000","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011100","101010001010","100101010101","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000100010","100001100111","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011010","011101000100","011100110011","100001010101","100001010101","100001010110","100101100110","100101100110","100101010110","011000110011","100001100111","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010101100","101010001001","011000110011","011101000100","011101000101","100001010101","100001010110","100101100110","100101100110","100101100110","011101000100","100001100111","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010101100","101010001010","011100110100","011101000100","011101000100","011101000100","100001010101","100001010110","100001010110","100101010110","011101000100","100101111000","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100110001010","101010011011","101010011011","101010101100","100110001001","100001010101","100001000101","011101000100","011101000100","011101000100","100001010110","011101000101","100001010101","100001010110","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100001010110","100001010101","100001010101","011101000101","011101000101","011101000100","100101100110","100101100110","100101010110","100101100111","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","100010001001","100110001010","101010011011","100101100111","100001000100","011101000101","011101000100","011101000100","011101000100","100001010110","100101100110","100101100110","100101100111","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011010","101010011011","100001111001","100001111001","100010001001","100001111001","100001100111","100001010101","011101000100","011101000100","100001010101","100101010110","100101100110","100101100111","100001111000","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100010001010","100110001010","101010011010","100110001010","100010001001","100110001001","100001010101","011101000100","011101000100","100001000101","100101010110","100101100110","100101111000","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011011","100010001001","100001111000","011101000101","011101000100","011101000100","100001010110","100101100110","100101100111","100101111001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","100110011011","100010001001","100001111001","100001100111","011101000100","011101000100","011101000100","011101000101","100001010110","100001100111","100001111001","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100110001001","100001100111","011101000100","011101000101","011101000101","100001010101","100101010110","100001100111","100110001001","100110001010","100001111000","100110001001","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100010001001","100110001010","100110001001","100001111000","100001100111","100101111000","100001100110","100001010101","011101000101","011101000101","100001010110","100001010110","100001100111","011001010101","100110001001","100110001001","100001111001","100110001010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010101100","100110011011","100110001001","100101111000","011101100111","011001000100","010100110011","010100110011","100001100110","011101010101","011001010101","011101000101","011101000101","100001010101","100001010110","100001111000","010000110011","010000110011","011001010101","100001100111","100101111001","100010001001","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100001100111","011101010101","010100110011","010000100010","001100100010","001100100010","010000100010","100001010110","011001010101","011001010101","100001010110","011101000100","011101000101","100001111000","011101100111","001100100010","001100100010","001100100010","001100100010","010101000100","011101100111","100001111000","100001111001"),
		("100110011011","100010001001","100110001010","011101100111","010000100010","001100100010","001100100001","001100100001","001100100010","001000100010","001100100010","100001100110","011001010101","011001010101","100001010110","011101000101","100001100111","100110001001","011101100111","001100100010","001100100010","001000100010","001000100010","001000100001","001000100010","010000110011","011101100111"),
		("101010011011","100110001010","100001111001","010101000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","011001000101","011001000101","011001010101","011101010110","100001111000","100110001001","100001111001","010000110100","001100100010","001100100010","001000100010","001000100010","001100100010","001100100010","001000100001","001100100010"),
		("101010101100","100110011010","100001111000","010000100010","001000100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001100110010","010101000100","011001010101","011001010101","011001010101","100001111000","011001010101","001100100010","001100100010","001000100010","001000100001","001100100010","011101000100","011101010101","010101000100","001100100010"),
		("100110011010","100110001010","100001100111","001100100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001","001100100001","001100100010","011001010101","011001010110","011001000101","011001010101","011001010101","010000110011","001000100010","001000100010","001000100010","001000100001","001100110011","100001010101","100001010110","100001010110","011001000100"),
		("100110001010","100001111001","011001000101","001100100010","001000100010","001100100010","001000100010","001000100001","001100100001","001100100001","001000100001","001100100010","011101100110","011101100110","010101000101","011001010101","010101000101","001100110011","001000100010","001000100010","001000100010","001000100001","010000110011","011101000101","100001010110","100001010110","011001000100"),
		("100110001010","100001111000","001100100010","001000100001","001000100001","001000100001","001100100001","001100100010","001000100010","001000100010","001000100010","001000100010","011101100111","011101100110","010101000101","010101000101","010101000100","001100100010","001000100010","001000100001","001000100001","001000100001","001100100010","011000110100","100001010101","100001010110","010100110011"),
		("101010011011","011101100111","001000100001","001000100001","001000100001","001000100001","001100100001","001000100010","001000100010","001000100001","001000100001","001000100001","011001010101","011001010101","010101000100","010101000101","010000110100","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","010100110011","100001000101","100001010101","010000110010"),
		("101010011011","011101100110","001000100001","001000100001","001000100001","001000100001","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","010000110011","010101000101","010101000100","010101000100","010000110011","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","010000110011","011101000101","100001010101","010000100010"),
		("101010011011","011001010101","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","001100100010","011101000100","100001000101","010000110011"),
		("100001111000","010101000100","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","001000100001","010000110011","010101000100","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","001000100001","001100100010","010000110011","001100100010"),
		("010101000100","001100100010","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","010100110011","011101000100","011001000100","011001000100","010101000100","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100100010","001100100010"),
		("001100100010","001100100001","001000100001","001000100001","001000010001","001000100001","001100100001","001000100001","010000110011","011101000100","011101000101","011101000100","011001000100","010000110011","010000110100","010000110011","001100100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001"),
		("001100100001","010000100010","001100100010","001100100001","001100100001","010000110011","001100100001","001100100001","011000110011","011101000100","011101000101","011101000101","011001000100","010000110011","010000110011","010000110011","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001"),
		("001100100001","001100100010","001000100001","001000100001","001100100010","001100100010","001000100001","001100100001","011000110011","011101000100","011101000100","011101000100","010100110100","010000110100","010000110011","001100110011","001000100010","001000100001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","001000010001","001000010001","000100010001"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000100010","010100110011","010000100010","001100100010","010000110011","010001000100","010000110011","001100100010","001000100010","001000100001","001000010001","001000010001","000100010001","001000010001","000100010000","000100010000","001000010001","001000010001","000100010000"),
		("001100100001","001000100001","001000100001","001000100001","001000100001","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001100110011","010000110100","010000110011","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","001000010001","001000010001","000100010000"),
		("010101000101","001100100010","001000100001","001000100001","001000100001","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010000110100","010000110011","001100100010","001000100001","001000010001","001000010001","000100010001","000100010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010000"),
		("101010011011","100110001010","011101100111","011001010101","011001010101","011001010110","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010000110011","010000110011","001100100010","001000100001","001000100001","000100010001","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000010001","001000010001"),
		("100110001010","100110011010","100110001010","100110001001","100101111000","100001100111","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001"),
		("100110001010","100110001010","100110001010","100110001001","100001111000","100001100111","001100100010","001000100001","001000010001","001000100001","001000100001","001000100001","001100110011","001100110011","001100100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001"),
		("100110001010","100110001010","100110001010","100110001001","100001111000","100001111000","010000110011","001000100001","001000100001","001000100001","001000100001","001000010001","001100110011","001100100010","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","000100010000","001000010001","001000010001","010101000100"),
		("100110001010","100110001010","100110001010","100110001001","100001111001","100001111000","001100110011","001000100001","001000100001","001000100001","001000100001","001000010001","001100110011","001100110011","001100100010","001000100010","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001100110011"),
		("100110001010","100110001010","100110001001","100110001001","100001111001","100001111000","001100110010","001000100001","001000100001","001000100001","001000010001","001000010001","001100110011","010101000100","010101000100","010000110011","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100001111001","100001111001","100001111000","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100110011","010001000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100001111001","100001111000","100001111000","100001111000","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100110011","010000110100","010101000101","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","100001111000","011101100111","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100110010","010000110011","010101000101","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010"),
		("011101100111","011101100111","100001100111","100001110111","100001111000","100001100111","001100110011","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","001100100010","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001"),
		("011101100110","011101100110","011101100110","011101100110","011101100110","011101100110","001100110011","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","001100100010","010000110100","010000110100","001100100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001"))
	-- 21
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100101111000","101010001001","100110001001","101010011010","101010011011","101010101100","101010011011","100110001010","100110001001","100110001001","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110001001","100101100101","100001000100","011101000011","011000110010","011000110011","100001010110","100110001001","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","100101111000","011000110010","010100100010","010100100010","010100100010","010100100010","010100100010","011101000100","100101111000","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010001001","100001010101","010100110010","010000100001","010000100001","010000100001","010000100010","010100100010","010100100010","011101010110","101010011011","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","100101111000","100001010100","011000110011","011000110100","011101000100","011101000100","100001010101","011101010101","011000110011","011001000101","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","101010011011","100101110111","011101000011","100001010101","100001010101","100101100110","100101100110","100101100110","100101100111","011101000101","011001000100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100110001010","101010101100","100001100111","011000110011","100001000101","011101000101","100001010101","100101100110","100101100110","100101100110","100001010101","011101000100","101010011010","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100110001010","100110001010","100101111001","011101000100","011101000100","011101000100","011101000100","100001010101","011101000101","100001010110","100001010101","011101010110","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","100010001001","100101111000","100001010101","011101000100","011101000100","011101000100","100001010110","100001010101","100001010110","100001010110","100001100111","100001111001","100110011010","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011010","101010011011","100001111001","100001010110","100101100110","100001000101","011101000100","011101000100","100001010110","100101100110","100101100110","100101100110","100101100111","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100010001010","100110001010","100101111000","100001010101","100001010101","011101000101","011101000100","100001010101","100101100110","100101100110","100101010110","100101111000","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","100101111001","100001010101","011101000101","011101000101","100001010110","100101100110","100101100110","100101111000","100110001010","100110001001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","100110011011","100110001001","100001010110","011101000101","011101000100","100001010110","100101100110","100101100110","100110001001","100010001001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100110001010","100110001010","101010011011","101010011011","100110001010","100001111001","100001010101","011101000100","011101000101","100001010110","100101010110","100001100110","100001111000","100001111000","100110001010","100110001010","100001111000","100110001001","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100001111001","100110001001","100110001010","100001111000","100101111000","100001010110","100001010101","011101010101","100001000101","100001010110","100001010110","100001111000","100110001001","101010011011","101010011011","100110001001","100001111001","100110001010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011100","100110001010","100010001001","100010001001","100001111001","100001111000","100001111000","100101100111","011101010101","011001010101","011001010101","100001010110","100001010110","100001010110","100001100111","100001111000","101010011011","101010011011","100110001010","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110001010","100110001001","100001111001","100001100111","011101010110","011101010101","100001100111","011101010110","011001010101","011001010101","100001010110","100001010110","100001010110","011101100110","010000110011","011001100110","100110001001","100110001010","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110001001","100001100111","011101000101","010100110011","001100100010","010000100010","100101111000","100001100111","010101000101","011001010101","100001010101","100001010101","100001100111","011001010110","001100100010","001100100010","001100100010","010001000100","011101100110","100101111000","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100001111000","100001100111","011001000100","010000110010","001100100010","001000100010","001000100001","001100100010","100101111000","100001100111","010101000101","011001010101","011101000101","011101010110","100110001001","011001010110","001100100010","001100100010","001100100010","001000100010","001000100010","010000110011","011001010110","100001111000","100001111001"),
		("101010011100","100001111001","010100110100","010000100010","001000100010","001100100010","001000100010","001000100010","001000100001","010000110011","100101111000","100001100111","011001010101","011001010101","100001100110","100101111001","100110001010","010101000101","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","010000110011","011101100111"),
		("100110011010","011101010110","001100100010","001100100010","001000100010","001100100010","001000100010","001000100010","001000100001","001100100010","011001000100","011001010110","011101100110","011101100110","100001110111","100110001001","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011"),
		("100010001001","011001000101","001000100010","001100100010","001000100010","001100100010","001000100010","001000100001","001100100001","001100100001","001100100001","010101000100","100001100111","011001010110","011001000101","011101010110","010000110100","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010"),
		("100110001001","010101000100","001000100010","001000100001","001000100001","001000100001","001100100001","001100100010","001000100010","001000100010","001000100010","010101000100","100001110111","011001010110","011001010101","010101000101","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001100100010"),
		("100110001001","010000110011","001000100001","001000100001","001000100001","001000100001","001100100001","001000100010","001000100010","001000100001","001000100001","010101000100","011101100110","011001010101","011001010101","010101000100","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001100100010"),
		("100110001001","001100100010","001000100001","001000100001","001000100001","001000100001","001100100010","001000100010","001000100001","001000100001","001000100001","010000110011","010101000101","011001010101","010101000101","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010"),
		("100001111001","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","011001000101","011001000101","010101000100","010000110011","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010"),
		("100001111000","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000101","010101000101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001100100010","011000110100","010101000100","001100100010","001000100001","001000100010","001000100010"),
		("100001111000","001100100010","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","011101000100","100001010110","011101010101","010000110011","001000100010","001000100010"),
		("100001100111","001100100010","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000010001","001100100010","010101000100","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","010000100010","100001000101","100001010110","100001010110","011001000100","001000100010","001000100010"),
		("100001100111","001100100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100010","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","010000110011","100001010101","100001010110","100001010110","010100110011","001000100010","001000100010"),
		("011001010101","001100100010","001000100001","001000100001","001000100001","001100100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","010000110011","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","001100100010","011101000100","100001010101","011101000100","001100100010","001000100001","001100100010"),
		("001100100010","001000100001","001000100001","001100100010","011001000100","011001000100","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010000110100","001100110011","001000100001","001000100010","001000100001","001000100001","000100010001","001000100001","011000110011","011101000100","010100110011","001000100001","001000100001","001000100010"),
		("010000110011","001100100010","011001000100","100001010110","100001010110","011000110011","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000100010","011000110011","010100110011","001000100001","001000100001","001000100010"),
		("010000110100","010100110011","011101000101","011101000100","011101000100","011000110100","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","000100010001","000100010000","000100010001","001000100001","001000100001","001000010001","001000100001","001000100010"),
		("010000110011","010100110011","011100110100","011000110011","011101000100","011000110100","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000100001","000100010001","000100010000","000100010000","000100010001","001000100001","001000010001","001000100010","001000100010","001000100001"),
		("001100100010","010000100010","011000110011","011100110011","011101000100","011000110100","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000100001","001100100010","001000100010"),
		("010101000100","001100100010","010000100010","011000110011","011000110011","001100100010","001000010001","001000100001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000010001","001000100001","001000100010"),
		("100110001001","011001010101","001100100010","010000100010","001100100010","000100010001","001000010001","001000100001","001000010001","001000010001","001000100001","001000010001","010000110011","001100110011","001000100010","001000100001","001000100001","001000100010","001000010001","000100010001","001000010001","001000010001","001000100001","000100010000","000100010001","001000010001","001100110011"),
		("100110001001","100110001001","011001010101","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","001100100010","001000100001","001000010001","001000100001","001000100010","001000100001","001000010001","001000100001","001000010001","010101000100","011001010101","010001000100","011001010101","100001111000"),
		("100110001010","100110001010","100001111000","001100100010","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","001000010001","010000110011","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000010001","010101000100","100110001001","100110001001","100110001001","100110001001"),
		("100110001010","100110001001","011101100111","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","010000110100","010101010101","010101000100","001100100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","010000110011","100101111000","100110001001","100110001001","100110001001"),
		("100110001001","100010001001","011001010110","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","010000110100","011001010101","010101000101","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100100010","011101100111","100110001001","100110001001","100110001001"),
		("100001111000","100001111000","011001010101","001000100001","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000110011","011001010101","010101000101","010000110011","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","010101000100","100001111001","100001111001","100001111001"),
		("011101100111","100001100111","010101000101","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","011001010101","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010001000100","100001111000","100001111000","100001111000"),
		("011101100110","011101100110","010000110100","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010101000100","010101000100","010000110011","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","010000110011","011101100111","011101100111","011101100111"))
	-- 22
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110011010","100110011011","100010001010","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010001010","101010001010","101010001001","100101111000","100110001001","100110011010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","100101111000","100101100101","100001010100","011100110011","011000110011","011101000100","100101100111","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001001","100001000100","011000110011","011000110010","010100100010","010100100010","011000110011","011000110011","100001010101","100110001001","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100101111000","011100110011","010000100001","010000100001","010100100010","010000100001","010100100010","010100100010","010100100010","100001100111","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100101110111","011101000011","011000110011","011000110011","011001000100","011101000100","100001010101","011101000100","010100100010","011101010101","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100101100111","100101010101","100001010101","100001010110","100101100110","100101100110","100101100110","100001010110","010100110011","011101010101","100110001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100101100111","100101010110","100001010101","100001010101","100001010110","100101100110","100101100110","100101010110","011000110011","011101010101","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011011","100110001001","100001010110","011101000100","011101000100","100001010101","011101000101","100001010101","100101010110","011100110100","100001010110","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100101111001","100001010101","011101000100","011101000100","100001010110","100001010101","100001010101","100001010110","011101000100","100001111000","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100101111000","100001010110","011101000101","011101000101","100001010110","100101100110","100101100110","100101100110","100001010110","100101100111","101010011011","100110001010","100110001001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100110001010","100110001010","100110001001","100001010110","011101000100","011101000100","100001010110","100101100110","100101100110","100101100110","100101100110","100101111000","100110011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100110001010","100110001010","101010011010","100101110111","011101000100","011101000100","100001010101","100101010110","100101100110","100101100110","100101111000","100110001010","100110001001","100001111000","100110001010","100110001010","100001111000","100110001010","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100010001001","100110001010","100101111001","011101000100","011101000100","100001010101","100001010110","100101100110","100101100110","100101111000","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100001111001","100110001010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011100","100110001010","100010001001","100010001001","100001111001","100001111000","100001010101","011101000100","011101010101","011101010101","011001010101","100001100110","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110001010","100001111001","100001111001","100101111001","100001111000","011101010101","011101000100","011101000101","011001010101","011001010101","100001100110","100001111000","100110001001","101010011010","100110011010","101010011011","101010011011","101010001010","100101111001","100001111000","100001111000","100001111000","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110001010","100001111001","100001111001","100110001001","100101111000","011101000100","011100110100","011101010101","011001010101","011001010101","100001010110","100001100111","011001010101","100001111000","100110001001","101010011011","101010011011","101010011010","100101111001","100101111001","100010001001","100001111000","100001111000"),
		("101010011011","100010001001","100001111001","101010011010","100110001010","100001111001","100001111000","011101010110","011101010110","011101000100","011101000100","011101000101","011001010101","011001010101","100001010110","100001100111","010000110011","001100100011","010000110100","011001010110","100001111000","100001111000","100001111001","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100001111001","100110001010","100110001001","100001010110","010100110011","001100100010","011001000100","100001100111","011101000100","011101000101","011001010101","011001010101","011101010110","100001111000","010000110011","001100100010","001100100010","001000100010","001000100010","001100110010","010101000101","100001100111","100110001001","100001111000","100001111000"),
		("100110001010","100010001001","100110001010","100001111000","011101000101","010000100010","001000100001","001000100001","010000110011","100101111000","100001100110","011101010101","011101100110","011101010101","100001100111","100110001001","010001000100","001100100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000100010","010101000100","100001111000","100001111000"),
		("100001111001","100001111000","011101010110","010100110011","001100100010","001000100010","001000100010","001000100001","010000110010","100001110111","100110001001","100001100111","100001100111","100001100111","100110001001","100001111001","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100001111001"),
		("011101100111","010100110100","001100100010","001000100001","001000100001","001000100001","001100100001","001100100010","001100100010","011101100110","011101100111","011101100111","100001111000","100001100111","100001111001","011001010110","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","011001010101","100001111001"),
		("010101000100","001100100010","001000100001","001000100001","001000100001","001000100001","001100100001","001000100010","001000100010","001100100010","010000110100","010101000100","011101010110","011001010101","010101000101","001100110011","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","010101000100","100101111001"),
		("010000110011","001100100010","001000100001","001000100001","001000100001","001000100001","001100100010","001000100010","001000100001","001000100001","010000110011","011001010101","011001000101","011001010101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010001000100","100110001001"),
		("010000110011","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100110010","010101000100","011001000101","010101000101","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","100101111001"),
		("010000100010","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","011001000101","010101000100","010000110100","010000110011","010100110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100001111000"),
		("001100100010","001100100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010101000100","010101000100","010101000100","010000110011","010000110011","011101000101","100001010110","011001000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000"),
		("001100100010","001100100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","010000110011","010101000100","010101000100","001100110011","010000110011","100001010101","100001010101","100001010110","010100110011","001000100001","001000100010","001000100010","001000100001","001000100010","001100100010","100001111000"),
		("010000110011","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001100110011","010101000100","010101000100","001100110011","010000110011","100001000101","100001010101","100001010101","010100110011","001000100010","001000100001","001000100001","001000100001","001000100001","001100100010","100001111000"),
		("010000110011","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001100100010","010101000100","010001000100","001100110011","010000100010","011101000100","011101000101","100001010101","010100110011","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","100001110111"),
		("010000110011","001100100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000010001","001100100010","010101000100","010101000100","001100110011","001000100001","001100100010","011101000100","011101010101","010100110011","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010101000100"),
		("100001010110","011101000100","001100100010","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","010001000100","010000110100","001100110011","001000100001","001000010001","010100110011","011101000100","010000110011","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010"),
		("100001010110","100001010101","011001000100","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110011","001100110011","001000100001","001000010001","001000010001","001100100001","001000100001","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010"),
		("100001010101","100001010110","100001010110","010000110010","000100010001","001000010001","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110100","010000110011","001000100001","001000010001","001000010001","000100010000","001000010001","001100100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100001"),
		("100001010101","100001010110","100001010110","011000110100","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110011","001100110011","001000100010","001000100001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001"),
		("011101000101","100001010110","100001010110","011001000100","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110011","010000110011","001100110011","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","001100100010"),
		("011000110100","100001000101","100001010101","010000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","010000110011","010000110011","001100110011","001000100010","001000100001","001000100010","001000010001","000100010001","001000010001","001000010001","000100010001","000100010001","000100010001","001000100001","011001010110"),
		("010100110011","010000100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","010000110011","010000110011","001100100010","001000100010","001000100001","001000100010","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001100100010","011001010110","100110001001"),
		("010000110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","010000110011","001100110011","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100001","010000110100","100001111000","100001100111","100001111000","100110001001","100110001001"),
		("011001010110","001100110011","010000110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001100110011","001100100010","001000100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100001","010000110011","100101111000","100110001001","100110001001","100110001001","100110001001"),
		("100001111001","100001111000","010101000101","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","010000110011","010101000100","010000110011","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001"),
		("100001111000","011101100111","001100100010","001000010001","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000110011","011001010110","011001010110","010101000101","010000110100","001100100010","001000100010","001000100001","001000100010","001000100010","011101100110","100110001001","100001111001","100001111001","100001111001"),
		("011101100111","011001010101","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","011001010101","011001010101","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100001","010101010101","100001111000","100001111000","100001111000","100001111000"),
		("011101100110","010101000100","001000010001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010101000101","010101000100","010101000100","010000110011","001100110011","001000100010","001000100010","001000100010","001000010001","010001000100","011101100111","011101100111","011101100111","011101100111"))
	-- 23
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010101100","101010101100","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","101010001001","101010001001","101010001001","101010001010","101010101100","101010011011","100110001010","100110001001","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","100101100110","100101010101","100001000100","011000110011","011101000011","100001100110","101010001010","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100101111000","011101000011","010100100010","010100100010","010100100010","010100100010","011000100010","011000110011","100001100111","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100101110111","011100110011","010000100001","010000100001","010000100001","010000100001","010100100010","010100100010","011000110011","100101111000","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100101111000","100001010101","011101000100","011000110011","011001000100","011001000100","011000110011","010100100010","010100100010","011101010110","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110001010","100101111000","100001010101","100001010101","100001010110","100101100110","100101100110","100101100110","011000110011","010000100010","011101010110","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100101100111","011101000101","100001010101","100001010110","100101100110","100101100110","100101100110","011000110011","010100100010","100001100111","101010011011","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100001010110","011101000100","011101000101","011101000101","100001010101","100101100110","100101100110","011000110011","010100110011","100101111000","101010011011","100110001010","100110001001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100110001011","100110001010","100001010110","011101000100","100001010101","100001010101","011101000100","100001010110","100101100110","011000110011","011001000100","101010001010","100110011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100110001010","100110001001","100001010101","100001000101","100101010110","100101100110","100001010110","100101100110","100101100110","011101000100","100001100111","101010011010","100110001001","100001111000","100110001010","100110001010","100001111000","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100001111001","100001010101","011101000100","100001010101","100001010110","100001010110","100001100110","100101100111","100001010110","100001100111","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100001111001","100110001010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011100","100110001010","100010001001","100101111001","100001010101","011101000100","100001010101","100001010110","100001010110","011001010101","011001010101","100001100110","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111000","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110001010","100001111001","100001111001","100001010110","011101000100","011101000101","100001010101","100001010101","011001010101","011001010101","100110001001","100110001001","100110001001","101010011010","100110011010","101010011011","101010011011","101010011010","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110001010","100001111001","100001111001","100001100111","011101000100","100001000101","100001010101","100001010101","011001000101","011101010110","100110001001","100001111001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011010","100101111001","100101111001","100010001001","100001111000","100001111000"),
		("101010011011","100010001001","100001111001","101010011011","100110001010","100001111001","100001111000","100001010101","011100110100","011100110100","011101000100","011101010101","010101000101","011001010101","100001111000","100001111000","100001111000","100001111000","100110001010","101010011011","101010011011","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001010","100010001001","100110001001","100101111000","011101010110","100001010110","011101000100","011100110011","011100110100","100001010101","100001010110","011001010101","011101100110","100001111000","100001111001","100001111001","100001111000","100001111001","100110001010","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("100110001010","100001111000","011101010110","010100110011","010000110010","010000100010","011101010110","011101010101","011100110100","011101000100","011101000101","100001010110","011101100110","100001100111","010101000101","011101100111","100110001001","100110001001","100001111001","100001111000","100001111000","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("011101010110","010100110011","001100100010","001100100001","001000100001","001000100010","011101010101","100001111000","011101000101","011101000100","011101000101","100001010110","100001100111","100001111000","010000110011","001100100010","010000110011","011101010110","100001111000","100001111001","100110001001","100001111001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001100100010","001000100010","001000100010","001000100001","001000100001","001100100010","100001100111","100110001001","100001100111","100001000101","100001000101","011101000101","100001111000","011101100111","001100100011","001100100010","001000100010","001000100010","001100110011","011001010101","100001111000","100110001001","100010001001","100001111001","100001111001","100001111001","100001111000"),
		("001000100001","001100100010","001000100001","001000100001","001000100001","001000100010","011101010110","100001111000","100001111000","100001100110","011101010110","100001111000","100001111000","011001010101","001100100010","001100100010","001100100010","001100100010","001000100001","001000010001","001100100010","011001010110","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001100100010","001000100001","001000100001","001000100001","001000100001","001100100010","010000110011","010101000100","011001010110","100001100111","100110001001","011101100111","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","011101100110","100110001001","100001111001","100001111000","100001111000"),
		("001000100010","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000101","010101000100","010101000100","011001010110","011001010110","001100100011","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000010001","010001000100","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","011001000101","011001010101","011001010101","011001010101","010101000101","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001100100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010101000100","011001010101","011001010101","011001010101","010101000100","001100110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100100010","100001111000","100010001001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110100","011001010101","011001010101","011001010101","010101000100","001100100011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100100010","100001111000","100110001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001100100001","001000100001","001000010001","001100100010","011001000100","011101000101","011101010101","011001010101","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001100100010","100001111000","100110001001","100110001001","100001111001"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010100110011","011101000101","100001010101","100001010101","011101010101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001100110010","100001111000","100110001001","100010001001","100101111001"),
		("001000100001","001000100001","001000100001","001000100001","001000010001","001100100010","011000110100","011101000101","100001000101","100001000101","011001000101","010001000100","010101000100","001100100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000010001","001100110011","100001111001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000100001","001000100001","000100010001","010000100010","011000110100","011101000100","011101000101","011101000100","010101000100","010000110100","010101000100","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100001","010000110011","100110001001","100110001001","100110001001","100110001001"),
		("001000010001","001000010001","001000010001","001000010001","000100010001","010000100010","011100110100","011000110011","010000100010","010000110011","010001000100","010000110100","010000110100","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100010","001000100001","010000110011","100110001001","100110001001","100001111000","100001100111"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","010000100010","010100100010","001100100001","000100010001","001000100001","010000110011","010101000100","010101000100","001100100011","001000100001","001000100001","001000100001","001000010001","000100010001","001000010001","001000100001","001000100010","001100100010","011101100111","100001110111","011001000100","011101000100"),
		("001000010001","001000010001","001000010001","001100100010","001000100010","001000100001","001000100001","001000010001","001000010001","001000100001","010000110011","010000110011","010001000100","001100110011","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","010000110011","011101000101","011000110011","011101000100"),
		("001000010001","001000010001","001000100001","001100100010","001000100001","001000010001","001000010001","001000100001","001000010001","001000100001","001100110011","010000110011","010000110100","001100110010","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000100010","011000110011","011000110100","011101010101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000100001","001100110011","010000110011","010001000100","010000110011","001000100001","001000010001","001000100001","001000100010","001000010001","000100010001","001000010001","001000010001","001000010001","010100100010","011000110011","011000110011","100001010101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","010000110011","010000110100","001100110011","001000100001","001000010001","001000100001","001000100010","001000100001","001000010001","001000100001","001000010001","001000010001","010100100010","011000110011","011000110011","011101000101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","010000110011","010000110011","001100110011","001000100001","001000010001","001000100001","001000100001","001000010001","000100010001","000100010001","000100010001","000100010000","001100100001","010000100010","010000100010","010100110011"),
		("010101000100","010101010101","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000100001","001000010001","001000100001","010000110011","010000110011","001100100011","001000100010","001000100001","001000100001","001000100001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","001000100001"),
		("100001111001","011101100111","001000100010","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001100100010","010000110011","001100100010","001100100010","001100100010","001000100001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000100001","010101000100"),
		("100001111000","011101100111","001000100010","001000100001","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000110011","001100110011","010000110011","010000110011","001000100010","001000100001","001000100001","000100010001","001000100001","001100110010","001100110010","001100110010","010001000100","011001100110","100001111000"),
		("011101100111","011101010110","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100100010","010001000100","010101000101","011001010101","010101000100","001100100010","001000100001","001000100001","000100010001","001000100001","011001010110","100001110111","100001111000","100001111000","100001111000","100001111000"),
		("011101100110","011001010101","001000100001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","001100100010","010101000100","010101000101","010101000101","010101000100","010000110011","001000100001","001000010001","000100010001","000100010001","001100100010","011001010110","011101100111","011101100111","011101100111","011101100111"))
	-- 24
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101110101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011011","101010011011","100110011010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010001010","101010011010","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001001","100101100110","100101010101","100001010101","100001010101","100101110111","101010011011","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001001","100001010101","011000110011","011000110011","011000100010","010100100010","011000100010","011101000100","100101111000","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011100","100110011011","100101110111","100001000100","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","100101111000","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110001011","100101100111","100001000100","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","100001100111","101010011010","100001111001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110001010","100001010101","100001010101","100001010101","100001010101","100001010101","100001010110","100101010110","011101000101","010100100010","100001100111","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101101","100110001001","100001010101","100001010101","100001010101","100001010101","100001010110","100101100110","100101100110","100101010110","011000110011","100001111000","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110001010","100101100110","100001010101","011101000100","100001010101","100001010101","100001010110","100101100110","100001010110","011000110011","100110001001","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100101111001","100101100111","100001000101","011101000100","011101000100","100001010101","011101000100","100001010101","100001010110","011101010101","101010011010","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100101111000","100101100110","100001010101","011101000100","100001010101","100101100110","100001010101","100101010110","100001010110","100001010110","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100101111001","100101100110","100001000101","011101000100","100001000101","100101010110","100101100110","100101100110","100101010110","100001100111","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100110001010","100110001010","101010101100","101110101100","101010011011","100110001010","100101111000","100001000101","011101000100","011101000101","100001010110","100001010110","100001100110","100101100110","100101111000","100010001001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011100","100110001010","100010001001","100101111001","100001010101","011101000100","011101000100","100001010101","100001010110","011001010101","011001010101","100101111001","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110001010","100010001001","100001111000","100001000101","011101000100","011101000101","100001010101","100001010101","011001010101","011001010101","100110001001","100110001001","100110001001","101010011010","100110011010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110001010","100001111000","100101100110","011101000100","011101000100","011101000100","100001010101","100001010101","011001010101","011001010101","100110001001","100001111001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011010","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100010001001","101010011010","100101111000","011101010101","100001010110","011101000100","011100110100","011000110011","100001000101","100001010101","010101000101","011001010101","100001111000","100001111000","100001111000","100001111000","100110001010","101010011011","101010011011","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","011101100111","011001000100","010100110011","010000100010","100001010110","011101000100","011100110011","011100110100","100001010101","100001010110","011001010101","011001010101","011001010110","100001111000","100001111001","100001111001","100001111001","100110001010","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("100001100110","010100110100","010000100010","001100100001","001100100001","001100100010","100001100111","100001100110","011100110100","011101000100","100001000101","100001010101","011101100110","011001010110","001100100010","001100110011","011001010101","100001111000","100001111001","100001111001","100001111000","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001100100010","001100100010","001000100010","001100100010","001000100001","001000100010","011101010110","100101111000","011101010101","011101000101","011101000101","011101010101","100001111000","011001010110","001100100010","001100100010","001000100010","001100110011","011001010101","100001111000","100110001001","100110001001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","011101100110","100110001001","100001111001","100001010110","100001010101","100001111000","100110001001","011001010101","001100100010","001100100010","001100100010","001000100010","001000100001","010000110011","011101100110","100001111001","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001100100010","001000100001","001000100001","001000100001","001000100001","010000110100","010101010101","011001010110","011101010110","100001110111","100110001001","100001111000","010101000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100001","001000100010","011101100110","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110010","011001010101","010101000101","010101000101","011101100111","011001010110","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","010101000100","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","011001010101","011001010101","011101010110","011001010110","011001010101","001100110011","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","010000110011","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010101000100","011001010101","011001010110","011001010110","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110100","011001010101","011001010101","011001010101","010101000100","001100100011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","100101111000","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","010000110011","011001010101","010101000101","011001010101","010101000100","001100100011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","100001111001","100110001001","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001100100010","010000100010","001000100001","001000100001","001000100001","001100100010","011001010101","010101000101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001100110011","100001111001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000100001","010100110011","100001010101","011000110011","001000100001","001000100010","001000100010","001100100010","011001010101","010101000100","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100001","001100100010","100001111000","100110001001","100110001001","100010001001","100101111001"),
		("001000100001","011001000100","011101000101","011101000100","011000110011","001100100010","001000100010","001000100010","001000100010","010101000100","010101000100","010000110100","010101000100","001100100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001100100010","100001111000","100110001001","100110001001","100110001001","100001111001"),
		("001100100010","011000110100","011000110011","011100110100","011001000100","001100100010","001000100010","001000100010","001000100010","010000110011","010101000100","010000110100","010101000100","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","011000110011","011000110011","011000110100","011000110100","001100100010","001000100010","001000100010","001000100001","001100100010","010101000100","010000110100","010000110100","001100100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100010","010000110011","100001110111","100110001001","100110001001","100101111001","100001111001"),
		("001000100001","010000100010","011000110011","011000110100","010100110011","001000100001","001000100001","001000100001","001000100001","001100100010","010000110100","010101000100","010000110100","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001000100010","010000110011","011000110100","011101100110","100101111001","100110001001","100010001001","100001111000"),
		("001000010001","001100100001","010100110011","011000110011","001100100001","001000010001","001000100001","001000100001","001000100001","001000100010","010000110011","010000110100","010001000100","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100100010","011000110011","011100110100","011101010101","100001111000","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001100100010","001100100010","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","010000110011","010000110100","010000110100","001100100010","001000010001","001000100001","001000100001","001000010001","001000010001","010000100010","011000110011","011101000100","011101000101","100001100111","100110001001","100110001001","100001111001"),
		("001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","010000110011","010000110011","010000110100","001100100010","001000010001","001000010001","001000100001","001000100001","001000010001","010000100010","011000110011","011101000101","100001010110","100001111000","100110001001","100110001001","100001111001"),
		("001100100010","001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","001100110011","010000110011","010000110011","001100100010","001000010001","001000010001","001000010001","001000010001","000100010001","010000100010","011000110011","011101000100","100001100111","100101111000","100110001001","100110001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001100100010","010000110011","010000110011","001100100010","001000100001","001000010001","000100010001","000100010000","000100010000","001000010001","010000100010","010100100010","011101010110","100110001001","100110001001","100110001001","100001111001"),
		("001000100001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000100001","001000100010","001100100010","010000110011","010000110011","001000100010","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","010101000101","100110001001","100110001001","100110001001","100001111001"),
		("001000100001","000100010000","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100010","001000100010","010000110011","010000110011","001100100010","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","001100100010","011101100111","100010001001","100110001001","100010001001","100010001001"),
		("001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","001100100010","010001000100","010101000100","010000110011","001100100010","000100010001","000100010000","001000100010","010101000100","010001000100","010101000101","011101100111","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100100010","011001010110","010101000100","010000110100","001100100010","001000010001","000100010000","001000010001","011001010101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000100010","010101000101","010001000100","010101000100","001100100010","001000010001","000100010000","000100010000","001100100010","011101100110","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 25
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100110001010","100010001001","100010001001","100110001011","100110011011","100110011011","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001001","100101111000","100101111000","100101111001","100001111001","100110001010","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110001010","100101110111","100101010101","011101000011","100001000100","011101000100","011101000100","100001010110","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101010101100","100101110111","100101010100","011000110010","010100100010","010100100010","010000100001","010100100010","010100100010","100001100111","100110011010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101010001001","100001010100","011000110010","010000100001","010000100001","010000100001","010000100001","010000100001","010100100010","100101110111","100110011010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","100110001010","011001000011","010100100010","010000100010","010000100001","010100100010","010100100010","010100110010","010100110011","011101000100","100110001001","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","100110001001","010100110010","010000100001","010000100001","010100110011","011101000100","100001010101","100101100110","100101100110","100101100110","100101111000","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101010011011","011000110011","010000100001","010100100010","011001000100","100001010101","100001010110","100101100110","100101100111","100101100111","100101111000","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101010011011","011000110011","010000100001","010100100010","011101000100","011101000101","100001010101","100001010110","100101100110","100101100110","100001100111","100110001001","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","101010011011","011000110011","010100100010","010100100010","011101000100","011101000101","011101000101","100001010101","100001010101","100101010110","100101100111","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110111101","101110101100","101010101100","101010101100","100001010110","011100110011","011000110011","011101000100","100001010101","100001010101","100001010110","100001010101","100001010110","100101111000","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110101101","100101111000","011101000100","011101000100","011101000100","011101000100","100001010101","100001010110","011101000100","100001010101","100101111000","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011011","101110101101","101010011011","100001010110","011101000100","011101000100","011101000100","011101000101","100001010101","100001010101","100001010110","100101111000","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100101111000","011101000101","011101000101","011101000100","011101000101","100001010101","100001010101","100101010110","100101111000","101010011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110001010","100101111001","100001000101","011101000100","011101000100","011101000100","100001010101","100001010110","100101100111","100001111000","100110001001","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","100110011011","100101111000","100001000101","011101000100","011101000100","011101000100","011101000100","100001010101","100001100111","100001111000","100001111000","100110001001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011011","100001100111","011001000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","011001010101","011001010101","011101100110","011101100111","100001111000","100110001010","101010011011","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100010001010","100010001001","100101111001","011101010110","010000100010","010000100010","011101010110","011101000100","011101000100","011101000100","100001010101","100001010101","011001010101","011001010101","010001000100","001100100010","010000110100","011001010110","100001111001","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110001001","011101100111","010100110011","001100100010","001000100001","001100100010","011101100110","011101010101","011101000100","011101000100","100001010101","011101000101","010101010101","011001010101","010001000100","001100100010","001100100010","001100100010","001100100010","011001010110","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("011001000100","010000100010","001000100010","001000100010","001000100010","001000100001","010101000101","100001111000","011101000101","100001010101","100001000101","011001000100","011001000101","011001010101","010000110100","001100100010","001100100010","001100100010","001100100010","001100100010","100001111000","100110001001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001100100010","001100100010","001000100001","010000110011","100001111000","100101111001","100001100110","011101000101","100001100111","011101100110","011001010101","001100110011","001100100010","001100100010","001100100010","001100100010","001100100010","011001010110","100001111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001100100001","001100100001","001000100010","001100110010","100001100111","100110001001","100001111000","011101100111","011101100111","011101100111","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010101000101","100110001001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001100100010","001100100010","001100100010","001100100010","001000100001","001000100010","001000100010","010101000101","011101100110","011001010110","011101100110","011001010101","011101100110","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010101000101","100110001001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001100100010","010101000101","011001010110","011001100110","010101010101","011101100111","011001010110","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","010101000100","100001111001","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","010101000100","011001010110","011001010110","010101000100","011001010101","010101000101","001100100010","001100100010","001100100010","001100100010","001000100010","001000100001","010001000100","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010000110011","011001010110","011001010101","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","011001010101","010101000101","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000101","010101000101","010001000100","010000110100","010101000100","010000110011","010000110011","001100100010","001000100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000100","010000110011","010000110011","010101000100","011101000100","011101010101","011101000101","001100100010","001000100010","001000100010","001000100010","100001100111","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100010","010000110011","010001000100","010000110011","001100110011","010100110100","011101000100","100001010101","100001010101","010000110011","001000100001","001000100010","001000100001","011001100110","100110001001","100110001001","100010001001","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001100110011","010001000100","001100110011","001100110011","010100110100","011101000100","100001010101","100001010101","010000110011","001000100001","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001100100010","010000110100","001100100010","001100100010","010000110011","011000110100","011101000101","011101010101","010000100010","001000100001","001000100010","001000100001","001000100001","011101100111","100110001001","100110001001","100010001001","100101111001"),
		("001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","001000100010","001000100010","001100100010","010000110011","001000100010","001100100010","001100100010","001000010001","010100110011","011101000100","001100100010","001000100001","001000100010","001000100001","001100100010","011101100111","100110001001","100110001001","100110001001","100001111001"),
		("000100010001","001000010001","000100010001","000100010001","000100010000","000100010000","000100010001","001000100001","001000100010","001100100010","010000110011","001000100001","001100100010","001100100010","000100010000","001100100010","010000100010","001000100001","001000100001","001000100001","001000100001","011001010110","100110001001","100110001001","100110001001","100110001001","100010001001"),
		("001000010001","000100010001","000100010001","000100010001","000100010001","000100010000","000100010000","001000010001","001000100001","001100100010","010000110011","001000100010","001100110011","001000100010","001000010001","001000100001","001000010001","001000100010","001000100010","001000010001","001100110011","100001111000","100110001001","100110001001","100110001001","100101111001","100001111000"),
		("001000010001","001000100001","010000100010","001100100010","001000010001","001000010001","000100010001","000100010001","001000010001","001000100010","001100110011","001000100010","001100110011","001100100010","000100010001","001000100001","001000100001","001000010001","001000100010","001100100010","011101100110","100110001001","100110001001","100101111001","100110001001","100010001001","100001111000"),
		("001000100001","010000100010","011000110100","011000110011","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","001100100010","001100110011","001100100010","001000010001","001000010001","001000100001","001100110010","011001010110","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("010100110011","011101000100","100001010101","011101000101","001100100010","000100010001","001000010001","001000010001","001000010001","001000100001","001100100010","001000100010","001100110011","001100100010","001000010001","001000010001","010000110011","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("010000100010","011000110011","011101000100","100001010101","010000100010","000100010001","001000010001","000100010001","001000010001","001000010001","001000100001","001000100001","001100110011","001100100010","001000100001","001000010001","001100110011","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100101111001","100110001001","100110001001","100001111001"),
		("001100100001","011000110011","011100110100","100001000101","010000100010","000100010001","001000010001","001000010001","001000010001","001000100001","001100100010","001100100010","001100110011","001100100010","001000100001","001000100001","001000100001","011101100111","100110001001","100110001001","100110001001","100110001001","100110001001","100101111001","100110001001","100110001001","100001111001"),
		("001000010001","001100100001","011000110011","011101000100","001100100010","000100010001","001000010001","000100010001","001000010001","001100110011","010101000101","010000110011","010000110011","001100100010","001000100001","001000100001","001000100001","010101000101","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000100001","000100010001","001000100001","001000100001","001000010001","001000010001","001000010001","000100010001","001000010001","010000110011","011001010101","010101000100","010000110011","001100100010","001000100001","001000100001","001000100001","010000110011","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000100001","000100010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","010000110011","011001010101","010101000100","010000110011","001100100010","001000100010","001000100010","001000100001","001100110011","100001111000","100110001001","100110001001","100110001001","100010001001","100010001001","100110001001","100010001001","100010001001"),
		("001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","010000110011","011001010101","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","011101100111","100010001001","100001111001","100001111001","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("000100010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010001000100","011001010101","010101000101","010000110100","001100100010","001000100001","001000100010","001000100010","001000100001","011001010101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010000","001000100010","001000100001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","010101000100","010101010101","010101000101","010000110011","010000110011","001000100010","001000100001","001000100001","001000010001","010001000100","011101100111","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 26
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100101111000","100101110111","100001100111","100001100111","100001111000","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100101111001","100101100110","100001000100","011000110011","010100100010","010100100010","010100110010","011000110011","100101111000","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110001010","100101100101","011101000011","010100100010","010000100001","010000100001","010000100001","010000100010","010100100001","011000110011","101010011010","101010101100","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001011","100110011011","100101100111","011101000011","010100100010","010000100001","010000100010","010000100001","010000100001","010000100001","010000100001","011000110011","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","100110001001","011001000011","010000100001","010000100001","010000100001","010100100010","011000110011","011000110011","011001000100","011000110011","100001100111","100110011010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","100001100111","010100100010","010000100001","010100100010","010000100001","011000110011","100001010101","100101100110","100101100111","100101100111","100101111000","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100001100110","010100100001","010000100001","010000100001","010100100010","011101000100","100001010101","100101100110","100101100111","100101100111","100101111000","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110011010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","100110001010","011101010101","010000100001","010000100001","010000100001","010100100010","011101000100","100001000101","100001010101","100001010101","100001010110","100101100111","101010011010","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","101010011011","011101010101","010100100001","011000110011","010100100010","010100110011","011101000101","100001010101","100001010101","100001010101","100001010101","100001100111","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101110101100","100001111000","011000110011","100001000101","011101000100","011100110100","011101000101","100001010101","100001010110","100101100110","100001010110","100001100111","100110001001","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","101010011010","011000110011","011101000100","011101000101","011101000100","011101000100","011101000101","100001010101","100101100110","100001010101","100001010110","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110111101","101010101100","101010101100","101010101100","100001100111","011100110011","011101000100","011101000100","011101000100","011101000101","100001010110","100001010110","100001010110","100101111000","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101010101100","101010011100","101010011011","101110101101","100110001001","011101000101","011101000100","011101000100","011101000100","011101000100","100001010101","100001010101","100001010101","100110001001","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011011","101010101100","101010011011","101010011010","100101111000","100001000101","011101000100","011101000100","011101000100","011101000100","011101000101","100001010101","100101100110","100110001001","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("100110001010","101010011011","100101111001","011001000101","100001010101","011101000100","011101000100","011101000101","011101000101","011101000100","011101000101","100001100110","100001100111","100001111000","100110011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100001111001","100001100111","010100110011","001100100001","011101010101","011101000101","011101000100","011101000101","011101000101","100001010101","100001100111","011101100111","100001100111","100001111000","100110001001","101010011011","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("010101000100","001100100010","001000100010","001000100010","011001000101","100001100110","011101000100","100001000101","100001010101","100001010101","100001100111","011001000101","011001010101","011101100111","011101100111","100001111000","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","100110011010","100010001001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","010000110011","100001111000","011101010101","100001000101","100001010110","011101000101","100001111000","011101100111","011001000101","011001010101","010101000100","001100100011","010101000101","100001111000","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100001","010000110010","100001111000","100001111001","100001010110","100001000101","011101000101","100110001001","100001111000","011001000101","011001010101","010101000100","001100100010","001100100010","001100110011","100001111000","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001100100010","001000100010","001100100010","011101100111","100110001010","100001111000","011101010110","100001111000","100110001010","011001010101","010101000101","011001010101","010101000100","001100100010","001100100010","001000100010","011001010110","101010011011","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001000100010","001000100010","010000110011","011001010110","011001010110","011101010110","011001100110","011001010110","010000110011","010101000100","011001010101","010101000100","001100100010","001100100010","001100100010","010101000100","100110001010","101010011010","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001100100010","001000100001","010001000100","011001010110","011001010101","011001010101","010101000100","001100100010","010000110011","011001010101","001100110011","001100100010","001100100010","001100100010","010000110011","100110001001","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001100100001","001100100001","001000100010","001100110011","011001010101","011001010110","011001010101","010101000100","001100100010","010101000100","011101100111","001100110011","001100100010","001100100010","001100100010","010000110011","100001111000","100001111000","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001100100010","001100100010","001000100001","001000100010","001100100010","010101000100","011001010101","011001010110","010101000100","001000100010","010101000101","100001100111","001100110011","001100100010","001100100010","001100100010","001100110011","100001111000","100110001001","100001111001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","010101000100","010101010101","011001010101","010001000100","001000100010","010101000101","100001110111","001100110011","001100100010","001100100010","001000100010","001100100010","100001111000","100010001001","100001111000","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010000110011","010101000101","010101000101","010000110100","001000100010","010000110011","010101000101","001100100010","001100100010","001100100010","001000100010","001100100010","100001111000","100001111001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000101","010101000100","010000110011","001000100010","001100100011","010000110011","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000100","001100110011","001000100010","001100110011","010000110011","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010000110100","001100110011","001000100010","001100110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100010","010000110011","011001000100","011000110100","010000110011","010000110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","010101000100","100101111000","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001100100010","010100110011","011101000100","011101000100","011101000100","011101000101","010000110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","010000110100","100101111001","100101111001","100110001001","100110001001","100010001001","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000010001","001000010001","001000100001","010100110011","011000110011","011101000100","011101000101","011101000101","011001000100","001100110011","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","010000110011","100101111000","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010100110011","011000110011","011101000100","011101000101","011101000101","010000110011","001100100010","010000110011","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000101","011101100111","011101010110","100001100111","100001111000","100101111001"),
		("001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","011000110011","011000110011","011101000100","011101000101","011101000100","001100100010","001100100010","001100110011","001000100001","001000100001","001000100001","001000100001","001000100010","001000010001","000100010001","001000010001","010000100010","011000110011","011101000100","011101000101","011101010110"),
		("000100010001","001000010001","000100010001","000100010000","000100010000","001000010001","010100100010","011000110011","010100110011","010100110011","010000100010","001000100001","001100100010","001100100010","001000100001","001000100001","001000010001","001000100001","001000010001","000100010000","000100010000","001000010001","010000100010","011000110011","011000110011","011000110011","011101000100"),
		("000100010001","000100010001","001000010001","001000010001","001000010001","000100010000","001000010001","001000010001","001000100001","001000010001","000100010001","001000100001","001100100010","001100100010","001000100001","001000100001","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","010000100010","011000110011","011000110011","011000110011","011101000100"),
		("001000010001","001000010001","001000010001","001100100010","001000100010","001000010001","000100010000","000100010001","001000010001","001000100001","001000010001","001000100001","001100100011","001100100010","001100100010","010000110011","001100100010","001000100001","000100010000","000100010000","000100010000","000100010000","001000010001","010100100010","011000110011","011000110011","011101000101"),
		("001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","000100010001","001000100001","001100110010","001100100010","001000010001","001000010001","011001010110","011101100111","010101000100","001100110010","001000100001","000100010001","000100010000","001000010001","001100100010","011001010101","100001111000"),
		("001000010001","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001100110010","001100100010","001000010001","001000010001","011001010101","100110001001","100110001001","100110001001","100001111000","011101100111","011001010110","010101010101","011001100110","100001111001","100010001001"),
		("001000010001","000100010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","001000100010","001000100001","001100110010","001100100010","001000010001","001000010001","010101000100","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001100100010","001000100001","001100110011","001100100010","001000010001","000100010001","001100110011","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100101111001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","001100110011","001000100001","001100110011","001100100010","001000010001","001000010001","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","010000110011","001000100010","001100100011","001100100010","001000100001","001000100001","001000100010","100001110111","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000010001","000100010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","001000100001","010000110011","001100100010","001100110011","001100100010","001000100010","001000100010","001000100001","011101100111","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001","100110001001","100010001001","100010001001"),
		("001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000100010","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001000100001","011001010110","100010001001","100001111001","100001111001","100001111001","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010101000100","010000110011","001100100010","001100100010","001000100001","001000100010","001000100001","010101000101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","000100010001","001000100010","010101000100","010000110011","001100100010","001000100010","001000100010","001000100001","001000100001","010000110011","011101100111","011101100111","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 27
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100010001001","100101111000","100101110111","100001100110","100001100110","100101110111","100001100111","100110001001","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110001011","100110001010","100101110111","100101010101","100001000100","011000110010","010100100001","010100100010","010100110010","011101000100","100101111000","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001010","100110011011","101010001001","100101100101","011000110011","010100100010","010000100010","010000100001","010000100001","010000100001","010100100010","011101000100","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010011010","100001010101","011000110010","010100100010","010000100001","010000100001","010000100001","010000100001","010000100001","010000100001","011101010101","101010011010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","100101111000","010100100010","010000100001","010000100001","010100100001","010100110010","011000110011","011001000100","011001000100","011101000100","100110001001","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100001010110","010100100001","010000100001","010000100001","010100100010","011101000100","100001010101","100101100110","100101100111","100101100111","100110001001","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110011010","100001111001","100001111001","100010001001"),
		("101110101100","101010101100","100110001010","011101010110","010000100001","010000100001","010000100001","011000110011","011101000101","100001010101","100101100110","100101100111","100101100111","100110001001","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","100110011010","011101010101","010000100001","010000100001","010000100010","011000110011","011101000101","100001000101","100001010101","100001010101","100001010110","100101100111","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101010101100","011101000101","010100100010","010100110010","010100100010","011000110100","011101000101","100001010101","100001010101","100001010110","100001010101","100001100111","100110001001","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","100101111000","011101000100","011101000100","011101000100","011101000100","011101000100","100001010101","100101010110","100101100110","100001010101","100101111000","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","101010011011","100001000101","011101000100","011101000100","011101000100","011101000100","011101000101","100001010110","100001010110","100001000101","100101111000","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101010101100","101010011100","101010011011","101110101100","100001100111","011101000100","011101000100","011101000100","011101000100","011101000100","100001010101","100001010110","100001010110","100110001001","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011011","101010011100","100110011011","101010101100","100110001001","011101000101","011101000100","011101000100","011101000100","011101000100","100001010101","100001010101","100001010110","100110001001","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("100110001010","101010011011","100110001010","100110001001","100101110111","011101000100","011101000100","011101000101","011101000101","011101000100","011101000101","100001010101","100001100111","100001111000","100110011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100010001001","100110001001","100101111000","011101000101","011101010101","011101000100","011101000100","011101000100","011101000101","011101000100","100001010101","100101111000","100101111001","100001111000","100110001001","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100001111000","011101100111","010100110011","001100100010","011101010101","011101000100","011101000100","011101000101","100001000101","100001010101","100001100111","100001111000","100001111000","100001111000","100001111000","100010001001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("010000110011","001100100010","001000100010","001000100001","011001010110","100001010110","011101000100","100001000101","100001010110","100001010101","100001100111","011001010110","011001000100","011001010101","011101100111","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100001","010101000100","100001111000","011101000101","100001010101","100001010110","011101000100","100001111000","011101100111","010101000101","011001010101","010101000100","010000110011","011101100110","100110001001","101010011010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001100100010","001000100001","010101000100","100001111001","100001111000","100001010110","100001000101","011101000101","100110001010","011101100111","010101000101","011001010101","010000110100","001100100010","001100100010","010000110011","100001111000","101010011010","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001000100010","010000110011","100001111001","100010001001","100001111000","100001010110","100001111000","100110001010","011001010101","010101000100","011001010101","010000110011","001100100010","001100100010","001000100010","010101000100","101010011010","101010011010","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","011001010110","011001010110","011001010110","011101100111","011101100111","001100100010","010001000100","010101000101","001100100011","001100100010","001100100010","001100100010","010000110011","100110001001","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001100100001","001100100001","001000100010","010101000101","011001010110","011001010101","011001010101","010101000100","001100100010","010101000101","011001010110","001100100010","001100100010","001100100010","001100100010","001100100011","100001111000","100001111000","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001100100010","001100100010","001000100001","001000100010","010000110100","011001010101","011001010110","011001010101","010000110100","001000100010","011001010110","011101100110","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100110001001","100001111001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","010000110011","010101000101","011001010101","011001010101","010000110011","001000100010","011001010110","011101010110","001100100010","001100100010","001100100010","001100100010","001000100010","011101100111","100110001001","100001111000","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010101010101","011001010101","010000110011","001000100010","010000110100","010101000100","001100100010","001100100010","001100100010","001100100010","001000100010","011101100110","100001111001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010001000100","010101000100","010101010101","010000110011","001000100010","001100110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000100","001100110011","001000100010","010000110011","010000110011","001000100010","001000100010","001000100010","001100100010","001000100010","011001010110","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010101000100","001100110011","001000100010","010000110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","010101010101","100110001001","100110001001","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110100","010000110011","001100100010","001000100010","010000110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100001","010001000100","100101111000","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001100110011","010000110011","001100100010","001000100010","001100110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100101111000","100101111001","100110001001","100110001001","100010001001","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000010001","001000010001","001000010001","001000100010","001100100010","010000110011","010101000100","010000110011","001000100010","001100110011","001100110011","001000100010","001000100010","001000100010","001000100001","001000100001","001100100010","100001111000","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","011000110100","011101000100","011101000101","011101000100","010000110011","001100110011","001100110011","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","100001100111","100110001001","100110001001","100110001001","100110001001","100010001001","100101111001"),
		("001000010001","001000010001","001000010001","001000010001","000100010000","010000100010","011000110011","011101000100","011101000101","011101000101","011101000100","001100100010","001100110010","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("000100010001","001000010001","000100010001","000100010000","000100010001","010100110011","011000110011","011101000100","011101000100","011101000100","010100110011","001000100001","001100110011","001100100010","001000100001","001000100001","001000010001","001000100001","001000010001","001000010001","010101000101","100001111000","100110001001","100101111001","100110001001","100110001001","100010001001"),
		("000100010001","000100010001","001000010001","001000010001","000100010001","010100100011","011000110011","011100110100","011101000100","011101000101","010000100010","001000100001","001100110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","000100010000","000100010000","001100100010","011001000100","011101000100","011101010110","100001010110","100001111000"),
		("001000010001","001000010001","000100010001","001000010001","001000010001","010000100010","011000110011","011000110011","011101000100","011000110011","001000100001","001000100001","001100110011","001100100010","001000010001","001000100001","001000010001","000100010001","000100010001","000100010000","000100010000","001000010001","010100100010","011000110011","011000110011","011000110011","011101000101"),
		("001000010001","000100010001","000100010001","001000010001","001000010001","001000100001","001100100001","001100100001","001100100010","001000100001","000100010001","001000010001","001100110011","001100100010","001000010001","001000010001","000100010001","000100010000","000100010001","000100010001","000100010001","001000100001","010100100010","011000110011","011000110011","011000110011","011101000100"),
		("001000010001","000100010000","001100100010","001100100010","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","000100010001","001000010001","001100110011","001100100010","001000010001","001000100001","001100100010","001000010001","000100010000","000100010000","000100010000","001000010001","010100100010","011000110011","011000110011","011000110011","011101000101"),
		("001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","001100100010","001100110011","001100100010","001000010001","001000010001","011001010101","011101100110","001100110010","000100010000","000100010000","000100010000","001100100001","010100100010","011000110011","011100110100","100001100110"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001100100011","001100110011","001100100010","001000010001","000100010001","010101000100","100110001001","100010001001","011001010110","001100110010","000100010001","000100010000","000100010001","011001000101","100001111000","100001111000"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","000100010000","001000100001","001100110011","010000110011","001100100010","001000010001","001000010001","001000100001","011101100111","100110001001","100110001001","100001111001","011101100111","010001000100","010000110011","100001111000","100110001001","100001111001"),
		("001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","010000110011","010000110011","001100100010","001000010001","001000010001","000100010000","011001010110","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000010001","000100010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","010000110011","010000110011","001000100010","001000010001","001000010001","001000010001","010101010101","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001","100110001001","100010001001","100010001001"),
		("001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","000100010001","001000010001","010000110011","010000110011","001100100010","001000100010","001000100001","001000010001","010101000100","100010001001","100001111001","100001111001","100001111001","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000100001","010000110011","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010000","001000010001","010000110011","010000110011","001000100010","001000100001","001000100001","001000100001","001100100010","011101100110","011101100111","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 28
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100010001001","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","100010001001","100110001010","100010001001","100010001001","100010001001","100001111001","100110001001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001010","100110011011","101010011011","100110001001","100101111000","100110001001","100101111000","100101111000","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010011011","101010011010","100101100110","100001010100","100001000100","011100110011","011100110011","011101010101","100101111000","100110001010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010011011","100101110111","011000110010","010100100010","010100100010","010100100010","010100100010","010100100010","011101000100","100110001001","101010011010","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100101111000","100101010101","010100110010","010000100001","010000100001","010000100001","010000100001","010100100010","010100100010","100001100110","101010011011","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101100","101010101100","100110001010","100001010110","011000110011","010100100010","010100100010","010100110011","011000110011","011101000100","011101000101","011000110011","011101000101","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","100110011011","100001100111","010100100010","011101000100","100001010101","100001010110","100101100110","100101100111","100101100111","100001010110","011101000100","100110001010","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101110101100","100001100111","011000110010","100001000101","100001010101","100001010101","100101100110","100101100110","100101100110","100101100110","011101000101","100101111000","100110001001","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","100101111000","011000110011","011101000101","011101000100","011101000100","100001010101","100001010110","100001010101","100001010110","100001100110","100101111001","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110101101","101010101100","101010011100","101010001010","011101000100","011101000100","011101000100","011101000100","011101000101","100001010101","100001010101","100001010101","100101100111","100110001010","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101010101100","101010011100","101010011011","100101111000","011101000100","011101000100","011101000100","011101000100","011101000100","100001010110","100101100110","100001010110","100101100111","100110001010","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011011","101010011100","101010011011","100110001001","100001000100","011101000100","011101000100","011101000100","011101000100","100001010101","100101100110","100001010110","100101111000","100110001001","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("100110001010","101010011011","100110001010","100110001010","100001100111","011101000101","011101000100","011101000101","011101000101","100001010110","100101100110","100001100110","100001111000","100001111000","100110011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100010001001","100110001001","100110001010","101010011010","100110001001","100001010110","011101000100","011101000101","011101000100","100001010101","100001010110","100101111000","100110001001","100001111000","100110001001","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100001111000","100001111001","101010011010","101010011011","100110001010","100001010110","011101000100","011101000100","011101000101","100001010110","100001010110","100101111000","100001111000","011101100111","100001111000","100001111001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100001111000","100001111001","100110001010","101010011010","100110001001","100001010101","011101000100","011101000100","011101000100","100001010101","100001010110","100001100111","011001010101","011001000101","011101100111","100001111001","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100001111001","100001111000","100110001001","100001111000","011001000100","011101010101","011101000100","011101000011","011101000100","100001000101","100001010110","100001100111","011001010101","011001010101","011101100110","011101100111","100001111000","100110001010","101010011010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110001010","100001111000","011001010101","010000100010","001100100010","011101010110","011101000100","011101000100","011101000100","011101000101","100001010101","100001100111","011001010110","011001010101","010101010101","001100100010","010000110011","010101010101","100001111000","101010011010","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("011101100110","010000110011","001000100010","001000100010","001000100010","011001100110","100001010110","011101000100","011101000101","011101000101","011101000100","100001111000","011001010110","010101000101","010101000101","001100100010","001100100010","001100100010","001100100010","010101000101","100110001001","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001100100010","001000100010","001000100010","001000100010","001000100010","010101010101","100110001001","011101010110","100001000101","011101000100","011101010101","100110001010","011101100111","011001010101","010000110011","001100100010","001100100010","001100100010","001100100010","001000100010","010101010101","100001111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001100100001","001000100001","010101000101","100010001001","100010001001","100001100111","011101010101","100001111000","100110001010","011001010101","011101100111","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","010000110011","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001100100010","001100100010","001000100001","010000110011","100001111000","100001111000","011101100111","011101100110","011101100111","011001010110","010000110100","100001100111","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100110011","100001111000","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100010","001000100001","001000100001","001000100010","001100110011","011001010101","011001010110","011001010101","011001010101","010000110100","010000110011","100001110111","001100110011","001100100010","001100100010","001100100010","001000100010","001000100010","001100100011","100001111000","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","010101000100","011001010110","011001010110","011001010101","010000110011","001100100010","010101000101","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","011001010101","011001010101","011001010101","010000110011","001100100010","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","011001010101","011001010101","010101000101","001100110011","001100100010","010000110100","001100100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010101000101","011001010101","010101000100","001100110011","001100100010","010000110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110100","010101000101","010000110100","001100100010","001100100010","010101000100","010100110011","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","011001010101","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010101000100","010000110011","001100100010","010100110100","011001000100","011101010101","100001010101","011101000101","001100100010","001000100010","001000100010","001000100001","010101010101","100110001001","100110001001","100010001001","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100001","001100100010","010000110011","010000110011","001100100010","011000110011","011001000100","011101000101","100001010101","100001010110","001100110011","001000100001","001000100010","001000100010","011001010110","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","001000100001","010000110011","010000110011","001100100010","010000110011","010101000100","011101000101","100001010101","100001010101","001100100010","001000100001","001000100001","001000100010","011101100111","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100001","001000010001","001000010001","001100110010","010000110011","001000100010","001000100001","010000110100","011000110100","100001000101","011101000101","001100100010","001000100001","001000100010","001000100001","001100110011","100001111000","100110001001","100110001001","100110001001","100001111001"),
		("000100010001","001000010001","000100010001","000100010001","000100010001","001000100001","001000100001","001000010001","000100010001","001100100010","010000110011","001000100010","001000100001","001100110011","001000010001","010100110011","010100110011","001000100010","001000100010","001000100001","001000100001","001000010001","011101100110","100110001001","100110001001","100110001001","100001111001"),
		("000100010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000100001","001000010001","000100010001","001000100001","010000110011","001000100010","001000100001","001100110010","000100010001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100001","010101000101","100101111001","100010001001","100001111001","100001111001","100101111000"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000100001","001100110011","001000100010","001000100010","001100100010","001000010001","001000100001","001000010001","001100100010","001000100010","001000100001","001100110011","100001111000","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000010001","000100010001","000100010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001100110011","001100100010","001100100010","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","011001010110","100110001001","100110001001","100110001001","100010001001","100010001001","100001111000"),
		("000100010001","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","001100100010","001100100010","001100110010","001000010001","001000010001","001000010001","001000100010","011001010101","100001111000","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001100100010","001100100010","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001100100010","001000100010","001100100010","001100110011","001000010001","001000010001","010001000100","100001110111","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001"),
		("011101000101","011101000101","001100100010","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","001000100001","001000010001","010000110011","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("011101000100","011101000101","010100110011","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","000100010001","001000100001","001000100010","010000110011","001100110011","001000100010","001000100010","001100100010","011101100111","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("011101000101","100001000101","011000110100","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","000100010001","001100110011","010101000100","010000110011","001100100010","001000100010","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("011101000100","100001000101","011001000100","001000100001","001000010001","001000010001","001000010001","000100010001","000100010001","000100010000","001100110010","010101000101","010101000100","010000110011","001000100010","001000100010","001000010001","001100110011","100001111001","100110001001","100110001001","100110001001","100010001001","100010001001","100110001001","100010001001","100010001001"),
		("011000110011","011101000100","011000110011","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","000100010000","001100100010","010101010101","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","011101100111","100010001001","100001111001","100001111001","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("001000100001","001100100001","001100100001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000100010","010101010101","010101000100","010000110011","001100100010","001000100010","001000100010","001000100001","010101010101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010000","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010000","001000100001","010101000100","010101000100","010000110011","001100100010","001000100001","001000100001","001000100001","010000110011","011101100111","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 29
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100010001001","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","100010001001","100110001010","100010001001","100001111001","100001111001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001010","100110011011","101010011011","100110001010","100110001010","100110001010","100010001001","100110001001","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010011011","101010101100","100110001010","100110001010","100110001010","101010011010","101010011011","101010011011","101010101100","101010011011","101010011010","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100110001010","101010011011","100101111000","100101100110","100001010101","100001010100","100001010101","100001100111","101010001001","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101100","101010101100","100110001010","101010011011","100101111000","100001000100","011101000011","011000110010","010100100010","010100100010","011000110011","011101000011","100001100110","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","101010011011","101010101100","100101110111","011000110010","010000100010","010100100010","010100100010","010000100001","010100100010","010100100010","011000110011","100101111000","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101010101100","101010101100","100101110111","011000110010","010100100010","010100100010","010100110011","011000110011","011101000100","011000110011","010100100010","100001010110","100110001010","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010011100","101010101100","101010101100","100101100111","100001000100","100001000101","100001010101","100101010110","100101100110","100101100110","100001010101","010100100010","011101010110","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110101101","101010101100","101010011011","101010101100","100001010101","100001010101","100001010101","100001010101","100001010110","100101010110","100101100110","100001010110","011000110011","011101010110","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101010101100","101010011100","101010011011","101010101100","100101100111","100001010101","011101000100","011101000101","100001010101","100001010101","100001010110","100001010110","011000110011","100001100111","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010101100","101010001001","100001010101","011000110011","011101000100","100001010101","011101000100","011101000101","100001010110","011101000100","100001111000","101010011011","101010011011","101010011011","101010011011","101010011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("100110011011","101010011011","100110001010","101010011010","100101111001","100001010101","011101000100","011101000101","100101010110","100101100110","100101100110","100101010110","100001010110","100001100111","100110011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100010001001","100110001001","101010011010","101010011010","100101100111","100001010101","011101000100","011101000100","100001010101","100101100110","100101100110","100101100110","100101100110","100001111000","100110001001","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100110001001","101010011010","101010011011","100110001001","100001010110","011101000100","011101000100","100001010101","100101100110","100001100110","100001010110","100001100110","100001111000","100001111000","100001111001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100001111000","100001111001","100110001010","101010011010","100110001010","100101100111","011101000100","011101000011","011101000100","100001010110","100001010110","100001010110","011001010101","011001010101","100001111000","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100001111001","100001111000","100110001001","101010011011","100110001010","100101111000","100001000101","011100110011","100001000101","100001010110","100001010110","011101010101","011001010101","011001010101","100110001001","100001111001","100001111001","100110001010","100110001010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110001010","100001111000","100110001001","101010011011","100110001010","100101111000","100001010101","011101000100","011101000100","100001000101","100001010110","011101010101","010101000101","011001010101","100110001001","100001111001","100001111001","100110001010","100110001010","101010011010","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("101010011010","100110001001","100001111001","101010011010","100110001001","100001111000","100001010101","011101000100","011100110100","011101000100","100001010101","011101010101","010101000100","011001010101","011001010110","011101100111","100001111000","100001111001","100110001010","101010011010","101010011010","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100001111001","100110001001","011101100110","011001000100","100001010101","011101000100","011100110011","011101000100","100001010110","100001010101","011001010101","010101000101","001100100010","001100100010","001100110011","010000110100","011001010101","011101100111","100001111001","100001111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("100110001001","100101111000","011101100111","010100110011","001100100001","010000110011","100001100111","011101000100","011101000100","011101000100","100001000101","011101000101","011101100111","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010000110011","010101010101","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100001100111","011001000100","001100100010","001000100001","001000100001","001100100010","100001111000","100001100110","011101000100","011101000101","011101000100","011101010110","100001111001","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","011001010101","100001111001","100010001001","100001111001","100001111000"),
		("010000110011","001000100010","001000100010","001000100001","001000100001","001100100010","011101100111","100010001001","100001100111","011101000101","011101000101","100001111000","100110001001","011001010101","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","010000110011","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100010","011101100110","100001111001","100001111000","011101010110","011101100111","100010001001","100001111000","010001000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000100","010101000100","010101000101","011001010110","011001010101","001100100011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101010101","011001010101","011001010101","011001010101","010101000101","001100110011","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","010101000101","100110001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","011001010101","011001010101","010101010101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010000110100","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010001000100","011001010101","011001010101","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100001111000","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","011001010101","010101010101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100010001001","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000100010","001000100001","001000100010","001000100001","001100100010","010101000101","010101000101","010001000100","010101000100","001100100011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","011101100111","100110001001","100001111001"),
		("001000100001","001000010001","001000010001","001000100001","001000100010","001000100001","001000100001","001000010001","001000100001","010101000100","010101000100","010001000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","011001010110","100110001001","100001111001"),
		("010100100010","001000010001","001000010001","001000010001","001000100010","001000100010","001000100001","001000010001","001000100001","010000110100","010101000100","010000110100","010001000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100001","011001010101","100110001001","100001111001"),
		("011101000100","010000100010","000100010001","000100010001","001000100001","001000100001","001000100001","001000010001","001000010001","001100110011","010101000100","010001000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001100100010","001000100010","001000100001","001100110011","011101100111","100010001001"),
		("100001010101","011000110100","001000100001","000100010001","001000010001","001000100001","001000100001","001000010001","001000010001","001100100010","010000110100","010000110100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","011000110011","010100110011","010000100010","001000100001","001100110011","100001111000"),
		("100001010110","100001000101","001100100010","000100010001","001000010001","001000100001","001000010001","001000010001","001000100001","001000100010","010000110011","010000110100","010000110100","001100100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001100100010","011000110100","011101000101","100001010101","010100110011","010101000100","100001111000"),
		("100001010101","100001010101","010000100010","000100010000","001000010001","001000010001","001000100001","001000010001","001000100001","001000100001","010000110011","010000110100","010000110100","001100110011","001000100001","001000100001","001000100010","001000100010","001000100001","001100100010","010100110011","011101000100","011101000101","100001010101","011101000101","011101100111","100001111001"),
		("100001010101","100001010110","010000100010","000100010000","001000010001","001000010001","001000010001","001000100001","001000010001","001000010001","001100110011","010000110011","010000110011","010000110011","001000100001","001000010001","001000100001","001000100001","001000100001","001100100001","010100110011","011101000100","011101000101","100001010101","100001010101","100001111000","100010001001"),
		("100001000101","011101000101","001100100001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","010000110011","010000110011","001000100001","001000010001","001000010001","001000010001","000100010000","000100010000","001100100001","010100110011","011101000100","100001010101","011101000101","100001100111","100110001001"),
		("010000100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010101000100","010000110100","010000110100","001100100010","001000100001","001000010001","000100010000","000100010000","000100010000","000100010000","001000100001","010100110011","011000110100","011001000100","100001111000","100010001001"),
		("001000010001","000100010001","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000010001","001000100001","010000110011","010000110100","010000110011","001100100010","001000100001","000100010001","001000010001","001000100001","000100010000","001000100001","001000010001","001000010001","001100100001","011001010110","100110001001","100001111001"),
		("001100100010","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","001100100010","010000110011","001100110011","001100100010","001000100001","001000010001","001000010001","001000100001","000100010000","010101000100","011001010110","001100110011","010101000101","100001111000","100110001001","100001111001"),
		("100001110111","011001010101","001000100001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010001","001000010001","000100010001","001100100010","010000110011","010000110011","001100110011","001000100010","001000100001","001000100001","001000100001","001000010001","010001000100","100110001001","100001111000","100001111000","100110001001","100010001001","100010001001"),
		("011101100111","001100110011","001000010001","000100010001","000100010001","001000010001","001000010001","000100010001","001000010001","000100010001","001000010001","010000110011","010101000100","010101000100","010101000100","010000110100","001000100010","001000100001","001000100001","001000100001","001100110011","100001111000","100001111001","100001111001","100001111001","100001111001","100001111001"),
		("011001010110","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000010001","010101000101","010101000101","011001010101","011001010110","010101000100","001100100010","001000010001","001000010001","001000100001","001000100010","011001010110","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("010000110011","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010000","000100010001","010001000100","010101000100","010101000101","010101010101","010101000100","010000110011","001000100001","001000010001","001000010001","001000100001","010101000101","011101100111","011101100111","011101100111","011101100111","011101100111"))
	-- 30
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100010001001","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","100010001001","100110001010","100010001001","100001111001","100001111001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001010","100110011011","101010011011","100110001010","100110001010","100110001010","100010001001","100110001001","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010011011","101010101100","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","101010101100","101010011011","101010011010","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100110001010","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","101010101100","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101100","101010101100","100110001010","101010011011","100110001010","100110001010","100110001010","100110011010","101010001001","100101110111","100101100111","100101100110","100101110111","101010001010","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","101010011011","101010101100","101010011011","100110001010","100110001010","100101110111","100001010100","100001000011","011000110010","010100100010","010100100010","011101000100","100101100111","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101110101100","101110101101","101010101100","100110001010","100110001010","100001010101","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","100001100111","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010011100","101010101100","101110101101","101010101100","100110001010","100101111000","100001000100","010100100010","010000100001","010100100010","010100110010","011000110011","011000110011","010100100010","011101000100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110111101","101010101100","101010011011","101110101100","101010101100","100110001010","100101111000","100001010100","011101000100","011101000101","100001010101","100001010110","100101100110","100101100110","011000110011","011001000100","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101100","101010101100","101010011011","101110101100","101010011100","100110001010","100001100111","100001000100","100001010101","100001010110","100001010110","100001010110","100101100110","100101100110","011101000101","011000110011","100110001010","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010101100","101010101100","101010011011","101010101100","101010011011","100110001010","100001100111","011101000100","100001000101","011101000101","100001010101","100001010101","100001010110","100101100110","100001010101","011001000100","101010011010","101010011011","101010011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","100110001010","101010011010","101010011011","100110001010","100101111000","100001010101","011101000100","011000110011","011101000101","100001010101","011101000100","100001010101","100001010101","011101010110","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100010001001","100110001010","101010011010","101010011010","100110001010","100110001010","100101111001","100101100111","011101000100","011101000100","011101000101","100101100110","100001010110","100101100110","100101010110","100001010110","100110001010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100110001001","101010011010","101010011011","100110011010","100110001010","100101111000","100101100110","100001000101","011101000100","011101000101","100001010110","100001100110","100001100111","100001100110","100001100110","100001111000","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100001111000","100010001001","101010011010","101010011010","100110001010","100110001001","100101111001","100101100111","100001010101","011101000100","011101000100","100001010110","011101010101","011001010101","011101010110","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110011010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100001111001","100001111000","100110001010","101010011011","100110001010","100101111001","100110001001","100110001001","100001010110","011101000100","011100110100","011101000101","011001010101","011001010101","100001111000","100001111001","100010001001","100110001010","100110001010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110001010","100001111000","100110001001","101010011011","100110001010","100001111000","100110001001","100110001010","100001100111","011101000100","011101000100","100001010101","011001010101","011001010101","100001111000","100001111001","100001111001","100110001010","100110001010","101010011010","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("101010011010","100110001001","100001111001","101010011010","100110001001","100001111001","100001111001","100110001001","100001100111","011101000100","011101000100","011101000101","011001000101","010101000101","100001110111","100001111001","100001111000","100001111001","100110001001","100110001010","101010011010","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100001111001","100110001010","100110001010","100001111001","100001111000","100110001001","100001010110","011100110011","011100110011","011101000100","011101010101","011001010110","100001100111","011101100111","100001111001","100001111001","100001111001","100110001010","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("100110001001","100101111001","100110001001","100110001001","100110001001","100001111000","100001100111","100001100111","100001010101","011101000100","011100110100","011101000101","100001100111","011101100111","100001100111","010101000100","010101000100","011101100111","100001111000","100010001001","100001111001","100110001001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100101111000","100101111000","100110001001","100001111000","100001100110","011001000100","010100110011","011101010101","100001010110","011101000100","011101000100","011101000100","100001100111","011101100111","100001100111","010101000101","001000100010","001100100010","010000110100","011001010110","100001111000","100110001001","100001111001","100001111000","100010001001","100001111001","100001111000"),
		("100110001001","100110001001","100001100110","011001000100","001100100010","001000100001","001000100001","011001000101","100101111000","011101000100","011101000100","011101000100","100001100111","100001111000","100001111001","010101000101","001000100010","001100100010","001000100010","001000100010","001100100010","010001000100","011101100111","100001111000","100010001001","100001111001","100001111000"),
		("100001100110","011001000100","001100100010","001000100001","001000100001","001000100001","001000100001","011001010101","100110001001","100001100111","011101000101","011101000100","011101010101","100001100111","100110001001","010001000100","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","010000110100","011101100111","100001111001","100001111000"),
		("001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","011001010101","100001111000","100010001001","100001100110","011101010101","011101100111","011101100111","100001110111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000101","011001010101","011101100111","011101100111","011101100110","010101000101","001000100010","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000100","010101000100","011001010101","010101000101","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100001111001"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000101","010101000101","010101000101","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100001111001"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000101","010101000101","010101000101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010101010101","100110001001"),
		("001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","010000110011","011001000100","010101000100","010101000100","010101000101","010101000101","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010000110100","100110001001"),
		("001000010001","001000010001","001000010001","001000100001","001100100010","011001000100","011101000101","011101000100","011000110011","010100110100","010101010101","010101000100","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100011","100001111000"),
		("001000100001","001000010001","000100010001","001000010001","011001000100","011101000100","011000110100","011000110100","010100110010","010000110011","011001010101","010101000100","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111"),
		("001000100001","001000010001","000100010001","001000100001","011101000100","011101000100","011101000100","011101000100","011101000101","011001000100","010101000101","010101000100","010101000100","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110"),
		("001000100001","001000010001","001000010001","001100100001","011000110100","011101000101","011101000101","011101000101","010100110011","001100100010","010001000100","010101000100","010001000100","010001000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","010001000100"),
		("001000100001","001000100001","001000100010","001100100010","011000110100","011101000101","011101000100","011001000100","001100100010","001000100001","001100110011","010000110100","010001000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001100100010"),
		("001100100010","001100100010","001000100001","001100100010","011000110011","010100110011","001100100001","001000010001","001000100001","001000100001","001100100011","010000110011","010001000100","010001000100","010000110011","001100100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010"),
		("001000100010","001000100010","001000100001","001100100001","010000100010","001100100001","000100010001","001000100001","001000100001","001000100001","001100100010","010000110011","010001000100","010000110100","010000110011","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001"),
		("001000100001","001000100010","001100100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","010000110100","010000110100","010000110011","001100100010","001000100001","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001"),
		("001000100001","001000100010","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","010000110011","010000110100","010000110011","001100110011","001000100001","001000010001","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001"),
		("001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000100001","001100100010","010000110011","010000110011","010000110100","010000110011","001100110011","001000100010","001000010001","001000100001","001000100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001"),
		("001000100001","001000100001","001000100001","001100100010","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","001000100010","010000110011","010000110011","010000110011","010000110011","010000110011","001000100010","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","000100010001","000100010001","001000010001","001000010001"),
		("011101100110","011001010110","011101100111","011101010110","001000010001","001000010001","001000010001","000100010000","001000010001","001000100001","001000100010","010000110011","010000110011","010000110011","010000110011","001100110011","001100100010","001000100001","001000100001","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010001","001000100001"),
		("100001111000","100001111000","100001111000","010101000101","001000010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001100100010","010000110011","010000110011","001100110011","010000110011","001100110011","001100100010","001000100010","001000100001","001000100001","000100010001","000100010000","000100010000","000100010000","001000010001","010000100010"),
		("100001110111","100001111000","100001111000","010000110011","000100010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001100100010","010000110011","010000110011","010101000100","010101000100","010000110011","001000100010","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000010001","010000100010"),
		("011101100111","011101100111","011101100110","001100100010","000100010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000100001","001100100010","010000110011","010101000100","010101010101","010101010101","010101010101","010000110100","001100100010","001000010001","001000010001","000100010001","000100010000","000100010001","001000100001","001000010001","010000100010"))
	-- 31

	);

	-- brick sprite
    type color_sprite is array (0 to 15, 0 to 15) of std_logic_vector(0 to 11);

    constant BRICK_ROM : color_sprite := (
        ("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
        ("000000000000","000100000000","001100000000","001100000000","001100000000","001100000000","001100000000","000000000000","001100000000","001100000000","001100000000","001100000000","001100000000","001100000000","001000000000","000000000000"),
        ("000000000000","001100000000","110000010000","101100010000","101100010000","101100010000","101000010000","001000000000","101000010000","101100010000","101100010000","101100010000","101100010000","101100010000","001100000000","000000000000"),
        ("000000000000","010000000000","110100010000","110100010000","110100010000","110100010000","101000010000","001000000000","101100010000","110100010000","110100010000","110100010000","110100010000","101100010000","001100000000","000000000000"),
        ("000000000000","010000000000","110100010000","110100010000","110100010000","110100010000","101000010000","001000000000","101100010000","110100010000","110100010000","110100010000","110100010000","101100010000","001100000000","000000000000"),
        ("000000000000","000100000000","001100000000","001100000000","001100000000","001100000000","001000000000","000000000000","001100000000","001100000000","001100000000","001100000000","001100000000","001100000000","000000000000","000000000000"),
        ("000000000000","001100000000","101100010000","100100010000","001000000000","011000000000","101100010000","101000010000","101000010000","101000010000","010100000000","001100000000","101100010000","100100010000","001000000000","000000000000"),
        ("000000000000","010000000000","111000010000","110000010000","001100000000","100000010000","111000010000","111000010000","111000010000","110100010000","011100000000","010000000000","111000010000","110000010000","001100000000","000000000000"),
        ("000000000000","001100000000","101100010000","100100010000","001000000000","011000000000","101100010000","101100010000","101100010000","101000010000","010100000000","001100000000","101100010000","100100010000","001000000000","000000000000"),
        ("000000000000","000100000000","001100000000","001100000000","001100000000","001100000000","001100000000","001000000000","000000000000","001100000000","001100000000","001100000000","001100000000","001000000000","000000000000","000000000000"),
        ("000000000000","010000000000","111000010000","110100010000","110100010000","110100010000","110100010000","100100010000","001000000000","110000010000","111000010000","110100010000","111000010000","110000010000","001100000000","000000000000"),
        ("000000000000","001000000000","011100010000","011100010000","100000010000","011100010000","011100010000","010100000000","000000000000","011100000000","100000010000","100000010000","011100010000","011000000000","001000000000","000000000000"),
        ("000000000000","000100000000","011000000000","010100000000","000100000000","001100000000","011000000000","011000000000","011000000000","010100000000","001000000000","000100000000","011000000000","010100000000","000100000000","000000000000"),
        ("000000000000","010000000000","111000010000","110000010000","001100000000","100100010000","111000010000","111000010000","111000010000","111000010000","011100000000","010000000000","111000010000","110000010000","001100000000","000000000000"),
        ("000000000000","001000000000","010000000000","010000000000","000100000000","001000000000","010000000000","010000000000","010000000000","010000000000","001000000000","000100000000","010000000000","010000000000","001000000000","000000000000"),
        ("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000")
    );

	-- apple gif sprite
	type apple_gif_sprite is array (0 to 1, 0 to 15, 0 to 15) of std_logic_vector(0 to 11);
	constant APPLE_GIF_ROM : apple_gif_sprite := (

		(	("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","000000000000","110010100010","000000000000","000000000000"),
		("000000000000","111111000011","111111000011","110010100010","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111111000011","111111000011","110010100010","000000000000"),
		("000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","100001010011","000000000000","000000000000","110010100010","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","100001010011","011001110011","000000000000","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","000000000000","111001110110","111001100110","000000000000","100001010011","011101000010","011001100011","011001110011","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","111001110111","111001100110","110100110011","110100110011","011101000010","010001100010","010001100010","110000110010","110000110011","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","111001110111","111001100110","111000110011","111110101010","111000110011","110000100010","110000100010","110000100010","111000110011","110100100010","110000110011","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","111001100110","111001000100","111110101010","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","110100100010","101100110011","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","111001010101","111000110011","111110101010","111000110011","111000110011","111000110011","111000110011","111000110011","110100100010","110000110011","101000110011","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","110100110011","111000110011","111110011001","111000110011","111000110011","111000110011","110100100010","110000110011","101000110011","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","110000110011","110100100010","111000110011","111000110011","111000110011","110100100010","110000110011","101000100010","100000100010","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","110010100010","000000000000","110000110011","101100110011","100100100010","000000000000","110000110011","101000110011","100000100010","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","111111000011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","110010100010","000000000000"),
		("000000000000","000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"))
	-- 0
	,

		(	("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111010110011","011101110000","000000000000"),
		("000000000000","000000000000","000000000000","111010110011","111101110000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111111110111","111111010100","111010110011","101110010010","000000000000"),
		("000000000000","111111110000","111111000011","111010110011","101110010010","000000000000","000000000000","000000000000","000000000000","000000000000","100101000011","111011001000","111111010101","111111000011","111111000011","000000000000"),
		("000000000000","111111010011","111010110011","110110100010","011101110000","000000000000","000000000000","000000000000","000000000000","100001010011","100001010011","100101100100","111111010101","111111010011","111101110000","000000000000"),
		("000000000000","111111110000","111010110011","000000000000","000000000000","111001100110","111001100110","000011111111","100001000011","100001010011","011001110011","010101110011","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","111001110111","111001100110","111001100110","110001000100","100001010011","011101000011","011001100011","011001100011","100101010011","111111110000","111010110011","111101110000"),
		("000000000000","111010110011","101101110011","111001110111","111001110111","111001100110","111001010101","110100110011","100001000011","010101100010","011001100010","110000110011","110000110011","110101100011","111010110011","101110010010"),
		("111111010100","111010110011","110110000100","111001110111","111001100110","111001100110","111010001000","111000110011","110100110011","110100110011","110100110011","111000110011","111000110011","110000110011","110101110010","000000000000"),
		("111111010101","111010110010","111001100110","111001100110","111001010101","111010011001","111001000100","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","101100110011","101100110011","111010110011"),
		("111111010100","111010110011","110101110100","111001010101","111001000100","111010011001","111001000100","111000110011","111000110011","111000110011","111000110011","110100110011","110000110011","101000100011","110110000011","111010110011"),
		("000000000000","111010110011","101101110011","110101010101","111000110011","111001000100","111001110111","111000110011","111000110011","111000110011","110100110011","110000110011","101000110011","101000100010","101101110011","111010110011"),
		("000000000000","000000000000","000000000000","101000100010","110000110011","111000110011","111000110011","110100110011","111000110011","110100110011","110000110011","101000100010","100100100010","011100100010","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","111100000000","110101010011","110000110011","110000100010","101000100010","110000110011","110000110011","101000110011","100000100010","100000100011","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","111111110000","111111000011","111010110011","110001100010","101100110011","100100100010","000000000000","110000100010","101000110011","100000100010","111111111111","111111010101","111111110011","111010110011"),
		("000000000000","000000000000","111111010011","111010110011","110110100010","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111111011001","111111010101","111111000010","111010110011"),
		("000000000000","000000000000","111111110111","111010110011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111111110111","111111010110","111111000011","111010110010"))
	-- 1

	);

	-- snale body sprite
	type color_sprite_8 is array (0 to 7, 0 to 7) of std_logic_vector(0 to 11);
	constant SNAKE_ROM : color_sprite_8 := (
		("010101100010","011010000010","011010000010","011010000010","011010000010","011010000010","011010000010","001001010001"),
		("011010000010","010011000001","001110110001","001110110001","001110110001","001110110001","001110110001","001001100001"),
		("011010000010","001110110001","000110100001","000110100000","000110100000","000110100001","000110100000","001001100001"),
		("011010000010","001110110001","000101110001","001010100001","001010100001","001001110001","001010100001","001001100001"),
		("011010000010","001110110001","000110100001","001010010001","001010010001","001010100001","001010110000","001001100001"),
		("011010000010","001110110001","000110100001","001010100001","001010100001","001010100001","001010110000","001001100001"),
		("011010000010","001110110001","000110110000","001010110000","001010110000","001010110000","001010110000","001001100001"),
		("001001010001","001001100001","001001100001","001001100001","001001100001","001001100001","001001100001","000101010001")
	);

--    vgaRed <= COLOR_ROM(row, col)(11 downto 8);

    constant img_size_x : natural := 16; -- size of the image sprites
    constant img_size_y : natural := 16;

    signal is_img_painted : std_logic;		-- is the rick gif painted
    signal img_clr : std_logic_vector(11 downto 0);

    signal img_x : unsigned(10 downto 0) := to_unsigned(50, 11); -- position of rick gif
    signal img_y : unsigned(10 downto 0) := to_unsigned(50, 11);
    
    signal rgb : std_logic_vector(11 downto 0); -- 12 bit rbg signal
    
    signal current_frame_gif : unsigned(11 downto 0) := to_unsigned(0, 12); -- the current gif frame from the array

    signal brick_clr : std_logic_vector(11 downto 0);  -- brick colour sognal

	signal snake_clr : std_logic_vector(11 downto 0); -- snake colour signal

	signal bcd_counter_out_1 : std_logic_vector(7 downto 0);  -- signals for the bcd counters
	signal bcd_counter_out_2 : std_logic_vector(7 downto 0);
	signal bcd_counter_1_cout : std_logic;
	signal bcd_counter_1_clk : std_logic;
	signal bcd_counter_2_clk : std_logic;
	signal increment_score : std_logic;
	signal bcd_counter_1_reset : std_logic;
	signal bcd_counter_2_reset : std_logic;

	signal is_gif_painted : std_logic;  -- is the gif painted
    signal gif_clr : std_logic_vector(11 downto 0); -- gif colour signal
	signal gif_x : unsigned(10 downto 0) := to_unsigned(212, 11);
    signal gif_y : unsigned(10 downto 0) := to_unsigned(50, 11);
begin
    led <= switch;  -- connect the leds to the switches
    start <= switch(7);
    
    process(pixel_clk) -- process to select the current frame of the GIF (can control the speed too)
    begin
        if rising_edge(pixel_clk)then
             if yCount = to_unsigned(1, yCount'length) and xCount = to_unsigned(1, xCount'length) then
                current_frame_gif <= current_frame_gif + 1;
             end if; 
        end if;
    end process;
    
	-- paint the apple gif at the current x, y position
    is_img_painted <= '1' when (xCount >= img_x and xCount < img_x + 16 and yCount >= img_y and yCount < img_y + 16) else '0';
    
	-- select the colours from the ROMs
	img_clr <= APPLE_GIF_ROM(to_integer(current_frame_gif(11 downto 3)), (to_integer(yCount - img_y) mod 16),(to_integer(xCount - img_x)) mod 16) when is_img_painted = '1' else (others => '0');

    brick_clr <= BRICK_ROM((to_integer(yCount) mod 16),(to_integer(xCount) mod 16)) when border = '1' else (others => '0');

	snake_clr <= SNAKE_ROM((to_integer(yCount) mod 8),(to_integer(xCount) mod 8)) when snakeBody /= (127 downto 0 => '0') else (others => '0');

	is_gif_painted <= '1' when (xCount >= gif_x and xCount < gif_x + 216 and yCount >= gif_y and yCount < gif_y + 384) else '0';
    gif_clr <= COLOR_GIF_ROM(to_integer(current_frame_gif(11 downto 3)), (to_integer(yCount(10 downto 3) - gif_y(10 downto 3)) mod 48),(to_integer(xCount(10 downto 3) - gif_x(10 downto 3))) mod 27) when is_gif_painted = '1' else (others => '0');

	-- instantiate BCD counter for minutes
    bcd_counter_unit_1 : entity work.nbit_bcd_counter(Behavioral)
        Port map (orig_clk => clk_100mhz, clk => bcd_counter_1_clk, up_down => '0', reset => bcd_counter_1_reset, cout => bcd_counter_1_cout, is_zero => open, output => bcd_counter_out_1);

    -- instantiate BCD counter for seconds
    bcd_counter_unit_2 : entity work.nbit_bcd_counter(Behavioral)
        Port map (orig_clk => clk_100mhz, clk => bcd_counter_2_clk, up_down => '0', reset => bcd_counter_2_reset, cout => open, is_zero => open, output => bcd_counter_out_2);

	-- instantiate four digits display
	four_digits_unit : entity work.four_digits(Behavioral)
		Port map (d3 => bcd_counter_out_2(7 downto 4),
                  d2 => bcd_counter_out_2(3 downto 0),
                  d1 => bcd_counter_out_1(7 downto 4),
                  d0 => bcd_counter_out_1(3 downto 0),
                  ck => clk_500hz, seg => seg, an => an, dp => dp);

	-- process to set the state of the bcd counters for the score
	process(clk_100mhz)
	begin
		if rising_edge(clk_100mhz) then
			bcd_counter_2_clk <= bcd_counter_1_cout;
			if game_over = '0' then
				bcd_counter_1_reset <= '0';
				bcd_counter_2_reset <= '0';
				if increment_score = '1' then
					bcd_counter_1_clk <= '1';
				else
					bcd_counter_1_clk <= '0';
				end if;
			elsif game_over = '1' then
				bcd_counter_1_clk <= '1';
				bcd_counter_2_clk <= '1';
				bcd_counter_1_reset <= '1';
				bcd_counter_2_reset <= '1';
			end if;
		end if;
	end process;

    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
        if pixel_clk = '1' then
            if start = '0' then -- intial start of the game conditions
                snakeX(0) <= to_unsigned(40, 7);
                snakeY(0) <= to_unsigned(30, 7);
                for count in 1 to 127 loop
                    snakeX(count) <= to_unsigned(127, 7);
                    snakeY(count) <= to_unsigned(127, 7);
                end loop;
                size <= to_unsigned(1, 7);
--                SIZE_INCREMENT <= 1;
                game_over <= '0';
            elsif game_over = '0' then
                if update = '1' then
                    for count in 1 to 127 loop
                        if size > count then
                            snakeX(count) <= snakeX(count-1); -- update the snake body position
                            snakeY(count) <= snakeY(count-1);
                        end if;
                    end loop;
                    case direction is
                        when "0001" =>
                            snakeY(0) <= snakeY(0) - to_unsigned(1, 7); -- update snake position based on the direction
                        when "0010" =>
                            snakeY(0) <= snakeY(0) + to_unsigned(1, 7);
                        when "0100" =>
                            snakeX(0) <= snakeX(0) - to_unsigned(1, 7);
                        when "1000" =>
                            snakeX(0) <= snakeX(0) + to_unsigned(1, 7);
                        when others =>
                            null;
                    end case;
                else 
                    if img_clr /= "000000000000" and (snakeBody /= (127 downto 0 => '0')) then                  
--                    if (snakeX(0) = pearX) and (snakeY(0) = pearY) then
                        img_x <= rand_X & "0000";  -- if food is eaten, increment size and change food position
                        img_y <= rand_Y & "0000";
                        if size < (128 - SIZE_INCREMENT) then
                            size <= size + SIZE_INCREMENT;
							-- double the size increment
--							SIZE_INCREMENT <= SIZE_INCREMENT * 2;
                        end if;
						increment_score <= '1';
                    
                    -- elsif border = '1' and snakeBody(0) = '1' then
                    elsif brick_clr /= "000000000000" and snakeBody(0) = '1' then -- border collision
                         game_over <= '1';
                    
                    elsif (snakeBody(127 downto 1) /= (127 downto 1 => '0') and snakeBody(0) = '1') then --snaek collision
                        game_over <= '1';

					else
						increment_score <= '0';
                    end if;
                end if;
            end if;
        end if;
        end if;
    end process;

	-- process to the direction of the snake based on the buttons
    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
            if pixel_clk = '1' then
            if (btn_up = '1' and direction /= "0010") then
                direction <= "0001";
            elsif (btn_down = '1' and direction /= "0001") then
                direction <= "0010";
            elsif (btn_left = '1' and  direction /= "1000") then
                direction <= "0100";
            elsif (btn_right  = '1' and direction /= "0100") then
                direction <= "1000";
            end if;
            end if;
        end if;
    end process;

	-- process to select level based on switch input
    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
        if pixel_clk = '1' then
            if switch(0) = '1' then
                if ((xCount(9 downto 3) = 0) or (xCount(9 downto 3) = 79) or (yCount(9 downto 3) = 0) or (yCount(9 downto 3) = 59) or ((xCount(9 downto 3) = 10) and (yCount(9 downto 3) >= 10 and yCount(9 downto 3) <= 20)) or ((xCount(9 downto 3) = 69) and (yCount(9 downto 3) >= 39 and yCount(9 downto 3) <= 49)) or ((yCount(9 downto 3) = 10) and (xCount(9 downto 3) >= 10 and xCount(9 downto 3) <= 20)) or ((yCount(9 downto 3) = 49) and (xCount(9 downto 3) >= 59 and xCount(9 downto 3) <= 69))) then
                    border <= '1';
                else 
                    border <= '0';
                end if;
            elsif switch(1) = '1' then
                if ((xCount(9 downto 3) = 0) or (xCount(9 downto 3) = 79) or (yCount(9 downto 3) = 0) or (yCount(9 downto 3) = 59) or((yCount(9 downto 3) = 20) and (xCount(9 downto 3) >= 10 and xCount(9 downto 3) <= 69)) or ((yCount(9 downto 3) =40 ) and (xCount(9 downto 3) >= 10 and xCount(9 downto 3) <= 69))) then
                    border <= '1';
                else 
                    border <= '0';
                end if;
            elsif switch(2) = '1' then
                if ((xCount(9 downto 3) = 0) or (xCount(9 downto 3) = 79) or (yCount(9 downto 3) = 0) or (yCount(9 downto 3) = 59) or ((xCount(9 downto 3) = 39) and (yCount(9 downto 3) >= 0 and yCount(9 downto 3) <=10)) or ((xCount(9 downto 3) = 39) and (yCount(9 downto 3) >= 49 and  yCount(9 downto 3)<=59))) then
                    border <= '1';
                else 
                    border <= '0';
                end if;
            else
                -- if (xCount(9 downto 3) = 0) or (xCount(9 downto 3) = 79) or (yCount(9 downto 3) = 0) or (yCount(9 downto 3) = 59) then
                if (xCount < img_size_x or xCount > 640 - img_size_x or yCount < img_size_y or yCount > 480 - img_size_y) then    
                    border <= '1';
                else 
                    border <= '0';
                end if;
            end if;
        end if;
        end if;
    end process;

	-- process to paint the snake body
    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
        if pixel_clk = '1' then
            for count in 0 to 127 loop
				-- change this to account for the size of the snake rom sprite which is 16x16
                if (xCount(9 downto 3) = snakeX(count)) and (yCount(9 downto 3) = snakeY(count)) then
                    snakeBody(count) <= '1';
                else
                    snakeBody(count) <= '0';
                end if;
            end loop;
        end if;
        end if;
    end process;
    
	-- set vgared, vgagreen, vgablue by splitting the 12 bit rgb signal
    vgared <= rgb(11 downto 8);
    vgagreen <= rgb(7 downto 4);
    vgablue <= rgb(3 downto 0);
    
	-- set the rgb signal based on the game state and the colours from the ROMs
    rgb <= (others => '0') when display = '1' else 
           gif_clr when game_over = '1' else
           snake_clr when (snakeBody /= (127 downto 0 => '0')) else
           brick_clr when border = '1' else 
           img_clr;

end Behavioral;