library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use ieee.math_real.all;
-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


entity snake is
    Port ( clk_100mhz : in STD_LOGIC;
           switch : in STD_LOGIC_VECTOR(7 downto 0);
           btn_up : in STD_LOGIC;
           btn_enter : in STD_LOGIC;
           btn_left : in STD_LOGIC;
           btn_right : in STD_LOGIC;
           btn_down : in STD_LOGIC;
           led : out STD_LOGIC_VECTOR(7 downto 0);
           vgared : out STD_LOGIC_VECTOR(3 downto 0);
           vgagreen : out STD_LOGIC_VECTOR(3 downto 0);
           vgablue : out STD_LOGIC_VECTOR(3 downto 0);
           hsync : out STD_LOGIC;
           vsync : out STD_LOGIC
         );
end snake;

architecture Behavioral of snake is
    signal pixel_clk : STD_LOGIC;

    constant SIZE_INCREMENT : integer := 4;
    
    signal xCount : unsigned(10 downto 0);
    signal yCount : unsigned(10 downto 0);
    signal rand_X : unsigned(6 downto 0);
    signal rand_Y : unsigned(6 downto 0);
    signal size : unsigned(6 downto 0);
    signal pearX : unsigned(6 downto 0) := "0101000";
    signal pearY : unsigned(6 downto 0) := "0001010";
    signal display : std_logic;
    signal R : std_logic;
    signal G : std_logic;
    signal B : std_logic;
    signal game_over : std_logic;
    signal pear, border : std_logic;

    type snake_array is array (0 to 127) of unsigned(6 downto 0);
    -- type snakeY_array is array (0 to 127) of unsigned(6 downto 0);

    signal snakeX : snake_array;
    signal snakeY : snake_array;

    signal snakeBody : unsigned(127 downto 0);
    signal update : std_logic;
    signal direction : std_logic_vector(3 downto 0);

    signal count : integer;

    signal start : std_logic;

    signal up, down, left, right : std_logic;

    signal grid : std_logic;

    type rom_type is array (0 to 15) of std_logic_vector(0 to 15);
    constant ROM : rom_type := 
    (
        "0000011111100000",
        "0001110101011000",
        "0010000010101100",
        "0110000000010110",
        "0100000001010110",
        "1000000000010011",
        "1000000000101111",
        "1000000000010101",
        "1000000001010011",
        "1010100001010111",
        "1010101010111011",
        "0101010101001010",
        "0111010111110110",
        "0011101101011100",
        "0001111011111000",
        "0000011111100000"
    );
    
    type color_gif_sprite is array (0 to 31, 0 to 47, 0 to 26) of std_logic_vector(0 to 11);
	constant COLOR_GIF_ROM : color_gif_sprite := (

		(	("100001111001","100001111001","100110001010","100001111001","100001111001","100010001010","100110011011","100110001010","100010001010","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100001111001","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100010001010","100010001010","100010001010","100010001010","100001111001","100001111001","100001111001","100010001010","100001111001","100001111001","100110001010","100110011011","100110011011","100110001010","100010001010","100010001010","100010001010","100010001010","100010001010","100010001010","100110001010","100110001010","100001111000","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100010001010","100010001010","100001111001","100001111001","100110011011","101010011011","101010101100","101010101100","101010011011","100110001010","100110001010","100110011011","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110011011","101010101100","101010011011","100110011011","100010001010","100010001010","100001111001","100110011011","101010011011","101010101100","101010101100","101010101100","101010101100","100110001010","100010001010","100010001010","100110001010","100110001010","100110011011","100010001010","100001111001","100001111001"),
		("101110101100","100110011011","100110001010","100110011011","100110011011","100110011011","101010101100","101010101100","100110011011","100110011011","100010001010","100110001010","101010011011","101010101100","101010101100","101010101100","101110101100","101110101100","101010011011","100110011011","100110001010","101010101100","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110001010","100110001010","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001010","100010001010","101010101100","101010101100","101010101100","101110101100","101110101100","101110101100","101010101100","100110011011","100110001010","101010011011","101010011011","100110001010","100010001010","100001111001","100001111001"),
		("100110001010","101010101100","100110011011","100110011011","100110011011","101010101100","100110001010","100010001010","100010001010","100010001010","100001111001","100010001010","100010001010","101010101100","101010101100","101110101100","101110101100","101010101100","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100110001010","100001111001"),
		("101010101100","101110101100","100110011011","100110011011","100110011011","100110011011","100110001010","101010101100","101110101100","101010101100","101010101100","100001111001","100010001010","101010011011","101010101100","101010101100","101010101100","101010011011","100110001010","100010001010","101010011011","101010011011","100010001010","100001111001","100001111001","100110001010","100001111001"),
		("101110101100","101110111101","100110011011","100110011011","100110011011","100110011011","101010011011","101110101100","101110101100","101010101100","101010101100","100110001010","100010001010","100010001010","100101100111","100001000011","100101100101","100101100111","100110001010","101010101100","101010101100","101010011011","101010011011","100010001010","100001111001","100001111001","100001111001"),
		("101110101100","101110111101","100110011011","100110011011","100110011011","101010101100","101110101100","101110101100","101010101100","101010101100","101010101100","100110001010","101010011010","100101100111","010100100010","010100100010","010100100010","011100110011","011000110011","101010011010","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("100110011011","101110101100","100110011011","100110011011","100110011011","100110011011","101110111101","101110111101","101110101100","101010011011","101010011011","100101111000","100101100101","100001000011","010100100010","010000100001","010000100001","010100100010","011000110011","011000110011","100110001001","100110011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","101110101100","101110101100","101110101100","101110101100","101010101100","101010011011","100101111000","100001000011","011100110011","010000100001","010000100010","010000100010","010000100001","010000100001","010000100001","011000110011","101010011010","100110011011","100110011011","100010001010","100001111001","100001111001"),
		("101110101100","100110011011","100110011011","100110011011","100110011011","101110101100","101110101100","101110101100","101110101100","101110101100","101010101100","100101100111","010100100010","011101000100","011101000100","100001010101","011000110011","010100100010","010100100010","010100100010","011000110011","101010011011","101010011011","100110011011","100110011011","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110011011","100110001010","100110011011","100110001010","101010101100","101010101100","101010011011","101010011010","100001000011","011000110100","100001000101","011101000101","100101100110","100101100110","100101100111","100101100111","011000110011","011000110100","101010011011","101010011011","100110011011","100110011011","100001111001","100001111001"),
		("101110101100","101110101100","100110001010","100110001010","100110011011","100110001010","100110001010","101010101100","101010101100","101010011011","100101111000","011100110011","011101000100","011100110011","011101000100","100101100110","100101100110","100101100110","100001010110","011101000101","100101111000","101010011011","101010011011","101010011010","100001111001","100001111001","100001111001"),
		("101110101100","101010101100","100110001010","100110001010","101010011011","101010101100","100110001010","100110001010","100010001010","100010001010","100001000101","100101100101","100001010101","011000110100","011000110100","011101000100","100001010110","100101100110","100001010110","011101000100","100110001001","101010101100","101010011011","100001111001","100001111001","100110001010","100001111001"),
		("101110101100","101010101100","100110001010","100110001010","100110011011","100110001010","100010001010","100010001010","100010001010","100001111001","100001000101","100101100101","100001010101","100001010110","100001010110","100001010101","100001010110","011000110100","100001010101","100001010110","100110001001","100010001010","100010001010","100001111001","100001111001","100110001010","100001111001"),
		("100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","101010011011","101010011011","101010011010","100010001010","100001010110","100101100101","100001010101","100101100110","011101000100","011101000101","100001010110","100001010110","100001010110","101010011010","100010001010","101010011010","101010011010","100001111001","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100010001010","100110001010","101010101100","101010011011","101010101100","100010001010","100101111000","100101100110","100001010101","011001010101","011001010101","011101000100","100001010110","100101100110","100101100110","101010011010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111000","100001111000"),
		("100001111001","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","100010001010","100001111000","100001111000","100001010110","100001010101","011101000101","011001010101","011001010101","100101100110","100001010110","100001010110","100101111000","100001111000","100010001010","100010001010","100110011011","100110011011","100110011011","100001111001","100001111000"),
		("100010001010","100001111001","100001111001","100001111000","100010001010","101010011011","101010011011","100110001001","100101111000","100101100111","011101000100","011101000100","011101000101","011001010101","011001010110","100001010110","100001010110","100010001010","100001111000","100001111000","100110001010","100110001001","100001111001","100110011011","100110011011","101010011010","100001111000"),
		("101010011011","100010001010","100001111001","100001111000","100001111000","101010011010","100110001010","100001111000","011000110100","100101100101","011100110011","011100110011","100001010110","010101000101","011001010110","100001010110","100101100111","100001111000","100001111000","100110001010","101010011010","100110001010","100001111001","100110001010","100110011011","100110001010","100001111001"),
		("101010011011","100110001010","100001111000","100001111000","100001100111","010100110011","010000100010","010000100010","010000100001","100001010110","011101000100","011101000100","011101000100","010101000101","011001010110","100001010110","100101111000","100001111000","100110001010","101010011010","101010011010","101010011010","100001111000","100001111000","100010001010","100001111000","100001111000"),
		("100110001001","011101010110","010100110100","010000100010","001100100001","001000100010","001000100001","001100100001","001100100001","100001100111","011101000100","011100110011","011101000100","011101100110","100001100111","100001010110","011101100110","100110001001","100110001010","100110001010","101010011010","101010011010","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("010000100010","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","100101111000","011101010110","011101000100","011101000100","100001111000","100101111000","100101111000","001100110011","001100110011","100110001001","100110001001","100110001010","100110001010","100110001010","100001111000","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010100110100","100001111000","100001111000","100001010110","100001000101","100101111000","100001100111","100110001001","001100110011","001100100010","001000100010","011101100110","100110001010","100110001010","100110001010","100001111000","100001111001","100110001001","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010101000101","100001111000","100110001001","100001010110","100001010110","011101010110","100001111000","100110001001","001100100010","001100100010","001000100010","001000100010","001100100010","100001111000","100001111000","100001111001","100110001001","100110001010","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001100110011","100001100111","100001111000","011001010110","100110001001","001100110011","001100100010","001000100010","001000100010","001100100010","001000100010","001100100010","100001111000","100001111000","100110001010","100110001010","100001111000"),
		("001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010110","010101000100","011001010110","011101100110","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010","001000100010","100001111000","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","011001010110","010101000100","010101000101","001000100010","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100010","100001111000","100001111001","100001111000","100001111000"),
		("001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100001111000","011001010110","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100001111000","100001111001","100110001001","100010001010"),
		("001000010001","001000010001","001000010001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","011001010110","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100101111000","100110001001","100001111001","100010001010"),
		("001100100001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","011101100110","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000010001","001000100010","001000100010","001000100010","100101111000","100110001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","010000110011","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100101111000","100010001010","100001111001","100001111001"),
		("001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","010000100010","010100110100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100110001001","100010001010","100010001010","100110001001"),
		("001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","010101000101","001100110011","010100110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100110001001","100110001001","100010001010","100110001001"),
		("001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","011001010110","001100110011","010100110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","100110001001","100010001010","100110001001","100001111001"),
		("001000100001","000100010000","001000010001","001000010001","001000010001","000100010000","001000010001","001000010001","001000100010","001000100010","001000100010","010101000101","010101000101","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","100110001001","100110001001","100110001001","100110001001"),
		("001000100010","001000010001","001000010001","001000010001","000100010000","000100010000","001000010001","001000010001","001000100010","001000100010","001000100010","011001010110","010101000101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001100100010","100110001001","100110001001","100110001001","100110001001"),
		("001000100010","001000010001","100001100111","100001010101","011101000100","010000100010","011000110100","011000110011","001000100010","001000100010","001000100010","011001010110","011001010110","010100110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","010000110011","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","011101000101","100101100111","100001010101","011101000100","011100110011","001100010001","001000100001","001000100010","001000100010","001000100010","010101000100","011001010110","010100110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","011101100110","100110001001","100110001001","100110001001","100110001001"),
		("001100100010","100101100111","100001010110","011101000100","011000110100","001100010001","000100010000","000100010000","001000100010","001000100010","001000100010","001000100010","010101000101","010100110100","001000100010","001000010001","001000100010","001000100010","001000010001","001000010001","001000100010","001000100010","100001111000","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","100101100111","100001010101","011100110011","001000010001","000100010000","000100010000","000100010000","001000100001","001000100001","001000100010","010101000100","010101000100","010100110100","001000100010","001000010001","001000100010","001000100010","001000010001","001000010001","001000010001","001000010001","001000100010","100110001001","100110001001","100110001001","100110001001"),
		("010000110011","100101100110","011000110100","001100010001","001000010001","000100010000","000100010000","000100010000","000100010000","001000100010","001000100010","001100100010","001100100010","010100110100","001000100010","001000010001","001000100010","001000010001","001000010001","000100010000","001000010001","001000100001","001100100010","100101111000","100110001001","100110001001","100110001001"),
		("001000100010","010000100010","001000100010","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000100010","001000010001","001000100001","010100110100","001100100010","001000100001","001000100001","001000010001","000100010000","001000010001","001000010001","001000010001","001100100010","100001111000","100110001001","100110001001","100110001001"),
		("001000100001","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000100001","001000010001","001000100010","010000110011","001100100010","001000100001","001000010001","001000100001","000100010000","000100010000","000100010000","001000010001","001000010001","011001010110","100001111000","100001111000","100001111000"),
		("001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","011001010110","011001010110","010100110100","001100110011","001000100010","001000010001","001000100001","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","010100110100","100001100111","100001111000"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","010101000101","010101000101","010000110011","001100100010","001000100001","000100010000","001000010001","000100010000","000100010000","000100010000","000100010000","001000010001","010000100010","011000110011","011000110011","011000110011"))
	-- 0
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100110001001","100110001010","101010011011","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100010001010","100001111001","100010001001","101010011011","101010011011","101010101100","101010101100","101010011011","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","100110001010","100010001010","100110001010","100110011011","101010011100","101010101100","101010101100","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010101100","101010011011","100110001010","100010001010","100110011011","101010011011","101010001001","100101110111","101010001001","101010011011","101110101100","101010101100","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100110001010","100010001010","100110001001","100101110111","011101000011","011100110011","011101000011","011101000100","100001100110","101010011010","101010011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110011011","101010011011","100110001010","100110001010","100110001010","100110001010","100001100111","100101100101","100001010100","010100100010","010000100001","010000100001","010100100010","010100100010","011101000100","100101111001","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001011","100110001011","100110011011","100110001010","101010011011","101010101100","101010011011","100001010101","011100110011","011000110010","010100100001","010000100001","010000100001","010000100001","010000100001","010100100010","100001100111","101010011011","100110011011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","100110011011","101010011011","101110101100","101110101101","101010011011","100001010101","010100100010","011000110011","011000110011","011000110011","010100110011","010100100010","010100100010","010100100010","100001100111","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010101100","101110101101","101110101100","101110101100","101010011011","011101000100","011000110011","011101000101","100001010101","100101010110","100101100110","100101100110","100101100110","011101000100","100001100111","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011100","101110101101","101110101101","101110101100","101010001001","011000110011","011000110011","011101000101","100001000101","100001010110","100101100110","100101100110","100101100111","100001000101","100001111000","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010101100","101110101101","101110101101","101010101100","100101100111","011100110011","011101000100","011101000100","011100110100","011101000100","100001010110","100101010110","100101100110","100001010101","100110001001","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101101","101010011100","100110011011","100110011011","100110011011","101010101100","101110101101","101110101101","101010011011","100001000101","011101000100","011101000101","011101000101","011101000101","011101000100","100001010101","011101000100","011101000100","100101111000","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110001011","100110011011","101010011011","101010101100","101010101100","100001010110","011101000101","011101000101","011101000101","100001010101","011101000101","100001010110","100101100110","100001100110","100101111001","100110011010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100110011011","100110011011","100110001010","101010011011","101010101100","101010001010","100001010110","011101000100","011101000100","011101000101","011101000100","100001010101","100101100110","100101100111","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010","100110001001","100001100110","011101000100","011101000101","011101000100","100001000101","100001010110","100101010110","100101111000","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100001111000","100001100111","011101000101","011101000100","100001000101","011101000100","100001000101","100001010101","100101100111","100110001010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100010001010","100110001010","101010011011","100001111000","011101000100","100001010101","011101000100","011101000100","100001010101","100001100110","100001100110","100001100111","100110001010","101010011010","100110011010","101010011010","100110001010","100110001010","100110011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110011010","100010001001","100010001001","100001111001","100001100111","011001010101","010000100010","010000100010","011101000101","011100110100","011101000100","011101010101","011001010101","011101010110","100110001001","101010011011","101010011010","100110001010","100110001010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100010001010","100110001001","100001101000","011101010101","010100110011","001100100001","001100100001","001000100001","001100100010","011001010101","011101000100","011101000100","011101010101","011001010101","011101100110","100110001001","101010011010","100110001010","100001111000","100001111001","100010001001","100110001010","100110011010","101010011011","100110011010","100010001001","100001111000"),
		("011101100111","011001000100","010000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","011001010110","100001100111","100001000101","011001010101","010101000101","011101100110","100001110111","010101000101","100001101000","100001111001","100010001001","100110001010","100010001001","100001111001","100110011010","101010011011","100110001010","100001111001"),
		("001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","100001111000","100001010110","011001000100","010101000101","100001100111","100001111000","001100100010","001100100010","010101000101","100110001001","101010011011","100110001010","100001111001","100110001010","100110011011","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","011101100111","100110001010","100001111000","100001010110","011001010101","100001111000","011101101000","001100100010","001100100010","001000100010","010000110011","011101101000","100110001010","100001111001","100001111001","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100001","001100100010","001100100001","011001010101","100001111001","100001111001","100001100111","100001111000","100110001001","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","011101101000","100110001001","100001111000","100001111000","100001111000","100001111001"),
		("001000100010","001100100010","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001100100010","011001010101","011001010110","011101100111","100001111000","100001111000","010000110011","001100100010","001100100010","001100100010","001100100010","001000100010","011001010110","100110001010","100001111001","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010","010101000101","011101100111","011101100111","100001111000","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010110","100110001010","100001111001","100001111001","100010001001","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","010101000100","011101100111","011101100110","011001010110","010101000101","001100100010","001100100010","001100100010","001000100010","001100100010","001000100010","010101010101","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010001000100","011101100111","011001010110","011001010101","010101000101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010101","100110001001","100001111001","100110001001","100110001010","100001111001"),
		("001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010000110011","011101100110","011001010110","011001010101","010101000100","001100100010","001100100010","001000100010","001100100010","001100100010","001000100010","011001010101","100110001001","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010000110011","011101100110","011001010110","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001100100010","001000100010","011001010110","100110001001","100001111001","100001111001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","011101100110","011001010110","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100010001001","100001111000","100001111001","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","011001010110","011001010110","010101000101","010001000100","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","011101110111","100010001001","100110001001","100010001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001100110011","011001010110","011001010101","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001100110011","100001111000","100110001001","100110001001","100010001001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100001","001100110011","011001010110","011001010101","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100010001010","100010001001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100001","001100110011","011001010101","010101000101","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100110001001","100010001010","100010001001","100110001001"),
		("001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001100110011","011001010101","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001"),
		("001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001100100011","010101000100","010101000100","010101000100","010000110011","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100010001001","100110001001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","001000100010","001100100010","010101000100","010101000100","010000110100","001100110011","001000100010","001000100010","001000100010","001000100001","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100110001001","100001111000"),
		("001000010001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","000100010001","001000100001","001000100010","001100100010","010000110100","010000110100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","011101100110","100110001001","100110001001","100110001001","100010001001"),
		("000100010000","000100010001","000100010001","000100010000","000100010000","000100010001","000100010000","000100010000","001000100001","001000100010","001000100010","010000110011","010000110011","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001100100010","011001010110","100010001001","100110001001","100110001001"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000100010","001000100010","001100110011","010000110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000010001","001000010001","011001100110","100110001001","100110001001"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","000100010001","001000010001","001000100001","001000100010","010000110011","010000110011","001100110011","001000100001","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000100001","000100010000","000100010000","001000100010","011001010101","100110001001"),
		("000100010001","000100010001","000100010001","000100010001","001000010001","001000010001","000100010000","000100010000","000100010001","001000010001","010000110100","011001010110","010101010101","010000110011","001000100001","001100100010","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","001000100001","010101000101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010001","001000010001","010101000101","011101100111","011001010110","010101000100","010001000100","010000110011","001100100010","001000010001","001000010001","010001000100","001100110011","001000010001","000100010001","000100010000","001000010001","010000100010","010100110011"),
		("000100010001","000100010000","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010101000101","011101100111","011001010101","011001010101","011001010110","010000110011","001000100010","001000010001","001000010001","011001010110","100001111000","010101000101","001000100001","000100010000","001000010001","010000100010","011000110011"),
		("001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010101000101","011101100111","011001010101","011001010101","011001010110","010000110100","001100100010","001000100001","001000010001","011001010110","100010001001","100001111001","011101100111","010000110011","001000100001","001000010001","010000100010"),
		("001000010001","001000010001","000100010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010101000101","011001100110","010101010101","011001010101","011001010110","010001000100","001100100010","001000010001","001000010001","011101100110","100001111000","100001111000","100001111000","100001111000","011001010110","001100110010","001000100001"),
		("000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000100001","010101000100","010101010101","010101000100","010101000100","010101010101","010000110100","001000100001","000100010001","001000100001","011001010110","011101100111","011101100111","011101100111","011101100111","011101100111","011101100110","011001010110"))
	-- 1
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001100110","100001010101","100101100110","100001100110","100101111000","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100101111001","100001100101","011000110010","011000110010","010100110010","010100100010","011000110010","011101010101","100110001001","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001001","100101100110","100001000011","010100100010","010000100001","010000100001","010100100010","010100100010","010100100010","100001100110","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011100","101010011011","100001010101","011100110011","011000110010","010100100010","010000100001","010000100001","010000100001","010000100010","010100100010","011101010101","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100001010101","010100100010","010100110010","011000110011","011101000100","011101000100","011101000100","011101010101","011101000100","011101000101","101010011011","101010011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110011011","101010011011","100110001010","100110001010","100001010101","010100100010","011101000100","100001000101","100001010101","100101100111","100101100111","100101100111","100101010110","011101010101","100110001001","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001011","100110001011","100110011011","100110001010","101010011011","100001010110","011000100010","011101000100","011101000101","100001010101","100001010110","100101100111","100101100111","100101010110","100001010110","100101111001","100110001001","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","100110011011","101010011011","101010101100","100001100110","011000110011","011101000100","011101000100","011101000100","011101000100","100001010101","100001000101","100001010101","100101110111","100110001001","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010101100","101110101101","101010011011","100001010101","011100110011","011101000100","011101000100","011101000101","011101000100","100001010101","100001010101","100001010110","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101101","101010011100","100001010110","011101000100","011101000100","011101000101","100001010101","011101000100","100001010101","100101100110","100101100111","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101010101100","101010101100","100101111001","100001000101","011101000100","011101000100","011101000100","011101000100","100001010101","100101100110","100101100111","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101101","101010011100","100110011011","100110011011","100110011011","101010101100","101110101100","101010101100","101010011011","100001100110","011101000100","011101000101","011101000100","011101000100","100001010110","100101010110","100101111000","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110001010","100110001010","101010011011","101010101100","100110001010","100001010110","011101000100","011101000101","011101000100","011101000100","100001010101","100101100110","100001111000","100001111000","100010001001","100110011010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100110011011","100110001010","100110001010","100001111000","011001000100","011101000101","011101000100","011101000100","011101000100","011101000101","100001010110","100101111001","100110001010","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","100110011011","100110001010","011101100110","010000110010","001100100010","011001000101","011101000100","011101000100","011101000100","011101000101","100001100111","100110001010","101010011010","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100001111000","011101010110","010100110011","001100100010","001100100010","001100100010","010101000101","100001010110","100001000101","100001010101","100001010101","100101100111","100110001010","101010011010","101010011010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110001001","011101010110","010100110011","001100100010","001000100010","001100100010","001100100010","001100100010","001100110011","100001111000","100001010110","100001010101","011101010110","100001100111","100001110111","011101100111","100110001010","101010011010","101010011010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("011001000101","010000110011","001100100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100001111000","011101010101","011001000101","011101100111","011101100111","001100100010","010000110100","100001111000","100110001010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("001100100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100001","001000100010","001000100010","011001010110","100110001010","011101010110","011001000101","100001100111","011101100111","001100100010","001100100010","001100110011","011101111000","100010001010","100110001010","100110001010","101010011011","100110011010","100010001001","100001111000"),
		("001000100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","001100100010","010000110011","100001111000","011001010101","010101000100","100001100111","011001010110","001100100010","001100100010","001100100010","011001010110","100110001010","100010001001","100001111001","100110011010","101010011011","100110001010","100001111001"),
		("001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010","010101000101","011001010101","011001010101","011101100111","010000110100","001100100010","001100100010","001100100010","011001010110","101010011011","100110001010","100001111001","100110001010","100110011011","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","010101000100","011001010110","011001010110","011001010110","001100110011","001100100010","001100100010","001000100010","011101100110","101010001010","100110001010","100001111001","100001111001","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001000100010","001100100010","001100100010","001000100001","001000100001","001000100001","001000100001","001100100010","001000100010","010000110011","011101100110","100001111000","011101100110","010000110011","001100100010","001100100010","001100100010","100001111000","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111001"),
		("001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001100100010","001100100010","001100110011","011101100110","100001111000","011101100110","010000110011","001100100010","001100100010","010000110011","100110001001","100110001001","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001100100010","001100100010","011001010110","100001111000","011101100110","010000110011","001100100010","001000100010","010101000100","100110001001","100110001010","100110001010","100110001010","100001111001","100001111001","100010001001","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001100100010","001100100010","010101000100","011101100110","011001100110","010000110011","001100100010","001000100010","010101000101","100110001010","100110001010","100110001001","100001111001","100001111001","100010001001","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","010000110100","011001010101","011001010110","010000110011","001100100010","001000100010","010000110100","100110001001","100110001010","100001111001","100001111001","100001111001","100110001001","100110001010","100001111001"),
		("001000100001","001000100001","001000100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","010000110011","011001010101","011001010110","010000110011","001000100010","001000100010","010000110100","100110001001","100001111001","100001111000","100010001001","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001100110011","011001010101","011001010101","010000110011","001000100010","001000100010","010000110100","100001111001","100001111001","100110001001","100110001001","100001111001","100001111001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","000100010001","001000010001","000100010001","000100010001","001000010001","001000100010","001100100010","010101000101","011001010101","010000110011","001000100010","001000100010","010001000100","100001111001","100110001001","100110001001","100001111001","100001111000","100001111001","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","000100010001","000100010001","000100010000","000100010000","001000010001","001000100010","001100100010","010101000101","010101000100","001100100010","001000100001","001000100010","010101000100","100001111001","100001111001","100001111001","100010001001","100110001001","100010001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010001","001000100001","001100100010","010101000101","010000110100","001000100001","001000100001","001000100010","010101000101","100001111001","100001111000","100001111000","100110001001","100110001001","100010001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001000010001","001100100010","010101000100","010000110011","001000100001","001000100001","001000100010","010000110011","100001111000","100001111001","100110001001","100110001001","100110001001","100010001010","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001100100010","010101000100","010000110011","001000100001","001000100001","001000100010","001000100010","010001000100","100001111000","100110001001","100110001001","100110001001","100010001010","100010001001","100110001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010001","001100100010","010000110100","010000110011","001000100010","001000100001","001000100010","001000100010","001000010001","010000110011","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001100100010","010000110100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000101","100001111000","100110001001","100110001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001100100010","010000110011","001000100001","001000100001","001000100010","001000100010","001000100001","001000100010","001000100010","001000010001","001100110011","100001111000","100110001001","100010001001","100010001001"),
		("001000100001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000100010","010000110100","001100100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000010001","001000010001","010101000100","100101111000","100101111001","100101111001"),
		("001000010001","000100010000","000100010001","000100010000","000100010000","000100010001","000100010000","000100010001","001000010001","000100010000","000100010000","000100010000","001000100001","010101000100","010000110100","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000010001","001100100010","011001000100","100001010101","100001010110","100001100110"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","001000100001","010101000100","011001010101","010000110100","001000100010","001000100010","001000100001","001100100010","001100110011","001000010001","001100100010","010100100011","011000110011","011000110011","011101000100"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","000100010001","001000010001","000100010000","000100010000","000100010000","001000100001","010101000100","011001010110","011001010110","001100110011","001000100010","001000010001","001100110011","100001111000","010101000101","001100100010","011000110100","011001000100","011000110011","011000110011"),
		("000100010001","000100010001","000100010001","000100010001","001000010001","001000010001","000100010000","000100010000","001000010001","000100010001","000100010000","000100010000","001000100001","010101000100","011001010110","011001010110","010001000100","001000100010","001000010001","001100100010","100001111000","100110001001","100001111000","100001111000","100101111001","100001100111","011101010101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001000100001","010000110100","011001010110","011101100110","010101000101","001000100001","000100010001","001100110011","100001111001","100110001001","100110001001","100110001001","100110001001","100110001001","100101111001"),
		("000100010001","000100010000","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001000100001","010000110100","011001010110","011101100110","010101010101","001000100001","000100010001","010001000100","100010001001","100010001001","100110001001","100110001001","100110001001","100110001001","100110001001"),
		("001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","000100010000","000100010000","001000100010","010101000100","011001010110","011101100110","010101000101","001000100001","000100010000","010101000101","100001111001","100001111001","100001111001","100001111001","100010001001","100010001001","100001111001"),
		("001000010001","001000010001","000100010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","000100010000","000100010000","001000100001","010101010101","011001010110","011001010110","010101000101","001000100001","000100010000","010101000101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000100001","010101000100","010101010101","011001010101","010101010101","001000100010","000100010001","010101000100","011101100111","011101100111","011101100111","011101100111","011101100111","011101100111","011101100111"))
	-- 2
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100001111001","100101111001","100101111000","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011010","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011100","100110001001","100101100110","100101100101","100001000100","011101000100","011101000100","100101100111","101010011011","101010101100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","100110001010","100101010101","011101000011","011000110010","010100100010","010100100010","010100100010","011000110011","100001100111","101010011011","101010011100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100101100111","011000110010","010000100001","010100100010","010100100010","010100100010","010000100010","010100100010","011001000100","101010011011","101010101100","101010011100","101010011011","100110011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110011011","100110001001","100101010101","011000110010","010000100001","010000100001","010000100001","010100110011","011101000100","011101010101","011000110011","100110001001","101010101100","101010011011","100110001001","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001011","100110011011","100101111000","011101000011","010100100010","011000110011","011101000100","100001010101","100001010110","100101100111","100101100111","011101000101","100001100111","101010011011","100110011010","100110001001","100110001001","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","100110001001","011000110011","011000110011","100001010101","100001010101","100101100110","100101100110","100101100111","100101010111","100001010110","100001111000","100110001010","100110001001","100110001001","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011011","011101000101","011000110011","011101000101","011101000101","100001010101","100001010110","100001010110","100001010101","100001010110","100101111000","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","100101111000","011000110011","011101000100","011101000100","011101000100","011101000101","100001010101","100001010101","100001010110","100101100111","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101010001010","011101000100","011101000100","011101000101","011101000100","011101000100","100101010110","100101100111","100101010110","100101100111","100110001010","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101101","101010011100","100110011011","100110011011","100110011011","101010101100","100110001001","011101000100","011101000100","011101000101","011101000101","011101000100","100001010101","100101100110","100101010110","100101111000","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110001010","100110001010","100110001010","100001010110","011101000100","011101000100","011101000101","011101000100","100001010110","100101010110","100101010110","100101111001","100001111001","100001111000","100010001001","100110011010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100110011010","100110001010","100110001010","100110001010","100001100111","011101000100","011101000100","011101000100","100001000101","100001010110","100101100110","100110001010","100110001010","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","100110011011","100110011010","100010001001","100110001001","100001100111","011101000100","011101000100","011101000100","100001010101","100101010110","100101100111","100110001010","101010011010","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100010001001","100001111001","100110001010","100110001001","100010001001","100001100111","011101000101","011101000100","011101000100","011101000100","011101000101","100001010101","100101100111","100110001010","101010011010","101010011010","100110011010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110001010","100001111001","100010001001","100010001001","100010001001","100110001001","010101000100","010000110011","011101000101","011101000100","011101000100","100001010110","100001100111","100001100111","100001111000","010101000101","011101100111","100110001010","101010011011","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100001111001","100001100111","010101000100","001100100010","001100100010","011101010110","100001010110","011101000101","011001010101","011001010101","011101010110","100001111000","010000110011","001100100010","010001000100","100001111000","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100001111001","100001111001","100101111000","011101010110","010000100010","001100100001","001100100001","001000100010","010000110100","100001111000","100001010110","011001010101","011001010101","011001010110","100001111001","010101000100","001100100010","001100100010","010000110100","100001111001","100110001010","100110001010","101010011011","100110011010","100010001001","100001111000"),
		("100001111001","100001111001","100001100111","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","011101100111","100001111000","011001000101","011001010101","011001010110","100110001001","010101000100","001100100010","001100100010","001100110011","100001111001","100010001001","100001111001","100110011010","101010011011","100110001010","100001111001"),
		("100101111001","011101010101","010000100011","001000100010","001000100010","001000100010","001100100010","001100100010","001000100010","001000100010","011001010110","100001111000","011001000101","011001010101","100001111000","100110001001","010000110100","001100100010","001100100010","010000110011","100110001010","100110001010","100001111001","100110001010","100110011011","100110001010","100001111001"),
		("010000110011","001100100010","001000100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001000100010","010000110011","100001111000","011101100110","011001010110","011101100111","011101100111","001100110011","001100100010","001000100010","010101000100","100110001010","100110001010","100001111001","100001111001","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","010101000101","011101100111","011101100111","011001010110","011001010110","001100110011","001100100010","001100100010","010101000101","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111001"),
		("001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","010000110011","100001100111","011101100111","011001010110","011001010110","010000110011","001100100010","001100100010","010101000101","100110001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100001100111","011001010110","011001010110","010000110100","001100100010","001000100010","010101010101","100110001010","100110001010","100110001010","100001111001","100001111001","100010001001","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001100100010","001100100010","001100100010","001100100010","010101000100","011101100110","011001010110","011001010110","010001000100","001100100010","001000100010","011001010110","100110001010","100110001001","100001111001","100001111001","100010001001","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","001000100010","001100100010","001100100010","001100100010","001000100010","010000110011","011001010110","011001010110","011001010110","010101000100","001000100010","001000100010","010101010101","100110001010","100001111001","100001111001","100001111001","100110001001","100110001010","100001111001"),
		("001000100001","001000100001","001000100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000100010","001100100010","001000100010","001000100010","010000110011","011001010110","011001010110","011001010110","010101000100","001000100010","001000100010","011001010110","100010001001","100001111000","100010001001","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100010","001100100010","001000100010","001000100010","010000110011","010101010101","011001010110","011001010110","010001000100","001000100010","001000100010","011001010110","100001111001","100110001001","100110001001","100001111001","100001111001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","010000110011","010000110011","011001010101","011001010101","010000110011","001000100010","001000100010","011101100111","100110001001","100110001001","100001111001","100001111000","100001111001","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","000100010001","000100010001","000100010000","001000100001","001000100010","001000100010","010000110011","001100110011","010101010101","011001010101","010000110011","001000100010","001100100010","011101100111","100110001001","100001111001","100010001001","100110001001","100010001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010001","001000100010","001000100010","010000110011","001100100011","010101000100","010101010101","001100110011","001000100010","001100100010","011101101000","100001111000","100001111000","100110001001","100110001001","100010001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000010001","001000100010","001100110011","001100100011","010000110011","010101000101","001100100010","001000100010","001100100010","100001111000","100001111001","100110001001","100110001001","100110001001","100010001010","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","001000010001","001100110011","001100110011","001100100011","010101000100","001100100010","001000100001","001000100010","011101010110","100110001001","100110001001","100110001001","100110001001","100010001010","100010001001","100110001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000010001","001100110011","001100100011","001100100010","010000110011","001000100010","001000100010","001000100001","001100100010","100101111000","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001100110010","001100100011","001000100010","001100100010","001000100001","001000100001","001000100010","001000100010","011001010101","100110001001","100110001001","100010001001","100110001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001100100010","001100100010","001000100001","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001100100010","001100100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","011001010110","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","000100010000","000100010001","000100010000","000100010000","000100010001","000100010000","000100010001","001000010001","001000010001","001000010001","000100010000","001100100010","001000100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100001","001000010001","010000110011","011101000101","100001100110","100001100111","100101111000","100110001001"),
		("001000100001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000100001","001000010001","000100010000","001100100010","001000100001","001000010001","001000100001","001000100001","001000100010","001000100001","001000100001","001000100001","010000100010","011000110011","011000110100","100001010101","100001010101","100001110111"),
		("001000100010","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","000100010001","001000010001","000100010000","000100010000","000100010001","001100100010","001000100001","000100010000","001000100001","001000100001","001000100001","001000100001","001000100001","000100010001","010000100010","010100100010","010100100010","011000110011","011101000100","011101000101"),
		("001100100010","000100010001","000100010001","000100010001","001000010001","001000010001","000100010000","000100010000","001000010001","000100010001","000100010000","000100010000","001100110010","001000100001","000100010000","001000010001","001000100010","001000100001","001000100010","011001010110","010000110011","011001010110","100001100111","011000110100","010100100010","011000110011","011101000100"),
		("001100100010","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","001000010001","000100010000","000100010000","001100100010","001000100001","000100010000","000100010000","001000100010","001000100001","001000100010","100001111000","100010001001","100110001001","100110001001","100001111000","011001000100","011101000100","100001100111"),
		("001100100010","000100010000","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001100100010","001000100001","000100010000","000100010000","001000100001","001000100001","001100110010","100001111000","100010001001","100010001001","100110001001","100110001001","100001111000","100001111001","100110001001"),
		("001000100010","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","000100010000","000100010000","000100010001","000100010000","000100010000","001100100010","001000100001","000100010000","000100010000","001000010001","001000010001","010001000100","100001111001","100001111000","100001111001","100001111001","100001111001","100010001001","100010001001","100001111001"),
		("001000100001","001000010001","000100010001","000100010001","000100010000","000100010001","001000010001","000100010001","000100010000","000100010000","001000010001","000100010001","001100100010","001000100001","000100010000","000100010000","001000010001","001000010001","010101000101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","001000100010","001000100001","000100010001","000100010000","001000100010","001000100010","010101000100","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111","011101100111","011101100111"))
	-- 3
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011010","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001001","100110001001","100110001001","100101111001","100001111001","100110001010","101010011011","101010011011","101010011100","101010101100","101010011100","101010011100","101010011011","100110011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001011","100101111001","100101110111","100101010101","100001010100","011101000100","100001010100","100001010101","100001100111","100110001001","101010011011","101010101100","101010101100","101010011100","101010011011","100110001001","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001001","100101010101","011101000011","011000110010","010100100010","010100100010","011000110011","011000110011","011000110100","100001111000","100110011010","101010011011","101010101100","101010011011","100110011010","100010001001","100110001001","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100001100110","011000110011","011000110010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","100001100110","100110001001","100110001010","101010011011","100110001010","100110001001","100110001001","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100001010110","010100100010","010000100001","010000100001","010100100010","011000110011","100001010101","100001010101","010100100010","011001000100","100110001001","100010001010","100110001001","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100101100111","011000110011","010100110010","011000110011","011101000101","100101010110","100101100111","100101100111","011101000100","011000110100","100110001010","100110001010","100110001010","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100101110111","011101000100","100001010101","100001010101","100001010110","100001010110","100101100111","100101100111","100001010110","011001000100","100110001001","100110001001","100110001001","100110001010","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100101111001","011101000100","011101000101","011101010101","100001010101","100001010101","100001010101","100001010110","100001010110","011101000101","100101100111","100001111001","100110001001","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110001010","100001010110","011101000100","011000110011","011101000100","100001010101","011101000101","100001010101","100101010110","100001010110","100101100111","100110001001","100110001001","100001111001","100001111000","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100101111001","100001010101","011000110100","011101000100","100001010110","100101010110","100101010111","100101010111","100101010110","100101100111","101010011010","101010011010","100110001010","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","100110001001","100001100110","011101000100","011101000100","100001010101","100001010111","100001010111","100101010111","100101100111","100110001001","100110011010","100110001010","101010011010","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001001","100110001010","100101100111","011101000101","011101000100","011101000101","100001010110","100001010110","100101010110","100101100111","101010011010","101010011011","101010011010","101010011010","100110011010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110001010","100010001001","100010001001","100010001001","100010001001","100001010110","011101000100","011101000100","100001010101","100001010110","100001010110","100001010110","100001111000","100110001010","101010011010","101010011010","101010011010","101010011010","101010011011","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100001111001","100110001010","100110001010","011101000101","011101000100","100001000101","100001010110","100001010110","011001010101","011001010101","011101100111","100001111000","011101100111","100001111000","100001111000","100110001001","100010001001","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100001111001","100001111000","100001111000","100110001001","101010011011","100110001001","011101010101","011101000100","011101000100","100001000101","100001010101","011001010101","011001010101","011101010110","001100100011","001100100010","001100100010","001100100010","010000110011","010000110100","011101101000","100110011010","101010011011","100110011010","100010001001","100001111000"),
		("100001111001","100001111000","100001111000","100001111000","100110001010","101010011010","011001000101","011001000100","011000110011","011000110011","011000110011","011101000101","011001010101","011001010101","100001111000","010000110100","001100100010","001100100010","001100100010","001100100010","001100100010","010000110100","100001111001","100110011010","101010011011","100110001010","100001111001"),
		("101010011011","100110001001","100001111000","100001111001","100110001001","011101010110","001100100010","011001000101","011101000100","011000110011","011100110100","011101000101","011001000101","011001010101","100001111000","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101101000","100110001010","100110011011","100110001010","100001111001"),
		("101010011011","100110001001","100001111001","100001111000","011001000101","001100100010","001000100010","010000110100","100001110111","011101010101","011101000100","100001000101","011001010101","011001010110","100110001001","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010110","100001111001","100010001001","100001111001","100001111000"),
		("101010011010","100110001001","100001100111","010100110100","001100100010","001100100010","001100100010","001100100010","011101100110","100001111000","100001100110","100001010110","011101010110","100001111000","100110001010","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010101","100001111001","100001111000","100001111000","100001111001"),
		("101010001010","100001100110","010000110011","001000100001","001000100001","001000100010","001000100010","001100100010","010101000101","100001111001","100010001010","100001111001","100001100111","100001111000","100110001001","010101010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011001010101","100001111001","100001111000","100001111000","100001111000"),
		("011001010101","001100100010","001000100001","001000100010","001000100010","001000100001","001000100010","001000100010","001100110011","011101100111","100001111001","011101100111","100001111000","100001100111","011101100111","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010101000101","100001111001","100001111001","100010001001","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010101","011001010110","011001010110","011101100110","011001010110","011001010101","001100110011","001100100010","001100100010","001100100010","001100100010","001100100010","010101000101","100001111001","100010001001","100110001010","100001111001"),
		("001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001000100010","010101000100","011001010110","011001010101","011001010101","011101100110","011001010110","001100110011","001000100010","001100100010","001100100010","001100100010","001100100010","011001010101","100010001001","100110001001","100110001010","100001111001"),
		("001000100001","001000100001","001000100010","001000100001","001000100010","001100100010","001100100010","001000100010","001000100010","001100100010","001100110011","011001010110","011001010101","011001010101","011001010110","011001010110","010000110011","001000100010","001100100010","001100100010","001100100010","001100100010","011101100111","100010001001","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","011001010101","011001010101","011001010110","011001010110","010000110100","001000100010","001100100010","001100100010","001100100010","001100100010","011101100111","100010001001","100001111001","100001111001","100001111001"),
		("001000100001","001000100001","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010101","011001010110","011001010110","011001010110","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100110011","100001111000","100010001001","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","010101000101","011001010110","011001010110","011001010110","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","100001111000","100010001001","100001111001","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010101","011001010110","011001010101","010000110100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","011101100111","100110001001","100001111001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000100010","001100100010","001000100010","001000100010","001000100010","001100110011","011001010101","011001010110","011001010101","010000110100","001100100010","001000100010","001100100010","001000100010","001000100010","001000100010","011001010110","100110001010","100010001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100001","001100110011","011001010101","011001010110","010101010101","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","010101000101","100110001010","100010001001","100110001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000100001","001000100010","001000100010","001000100001","001100110011","010101000101","011001010101","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","011101100111","100110001010","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010001","001000100001","001000100010","001000100010","001100110011","010000110011","011001010101","010101000100","010000110100","001100110011","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","010000110011","100001111000","100010001001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010000","001000010001","001000100010","001000100010","001100110011","001100110011","010101000100","010101000100","010000110011","001100100010","001000100001","001000100010","001000100010","001000100001","001000010001","001000010001","001000100010","100001111000","100110001001"),
		("001000100001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","001000010001","001000100010","001100110011","001100100010","010001000100","010101000100","010000110100","001100100010","001000100001","001000100001","001000100010","001000100001","000100010001","001000100001","001100100010","011101100111","100110001001"),
		("001000010001","000100010000","000100010001","000100010000","000100010000","000100010001","000100010000","000100010001","001000010001","000100010000","001000010001","001000100001","001100110011","001100100010","010000110011","010101000100","010000110100","001100100010","001000100001","001000100001","001000100010","001000010001","000100010000","001100100010","011001000100","011101000101","100001010110"),
		("001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001100110011","001100100011","001100100010","010000110100","010000110011","001100100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100001","011000110100","011000110100","011000110011"),
		("001000010001","000100010000","000100010000","000100010000","000100010000","001000010001","000100010001","000100010001","001000010001","000100010000","000100010000","000100010001","001100100010","001100100010","001000100010","010000110011","010000110011","001100100010","001000010001","001000100001","001000100001","001100110010","011101100110","001100100010","010000100010","011101000100","011101000100"),
		("001000010001","000100010001","000100010001","000100010001","001000010001","001000010001","000100010000","000100010000","001000010001","000100010001","000100010000","000100010000","001100100010","001100100010","001000100010","001000100001","001100100010","001100100010","001000010001","001000100001","001000100001","001100100010","100001111000","100001100111","010000100010","011000110011","100001010110"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","001000010001","000100010000","000100010000","001100100010","001100100010","001000100001","001000100010","010001000100","010000110100","001000100001","001000010001","001000100001","001100100010","100001111000","100110001001","011101010110","011001000100","011101010110"),
		("001000010001","000100010000","001000010001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001100100010","001000100001","001000010001","001100110011","011001010101","010101010101","010000110011","001000100010","001000100001","001000100010","011101110111","100110001001","100110001001","100001111000","100001111000"),
		("001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","000100010001","000100010000","000100010001","000100010000","000100010000","001100100010","001000100001","000100010000","001100100010","011001010101","011001010110","010101000101","001100110011","001000010001","001000100010","011101100111","100010001001","100010001001","100010001001","100010001001"),
		("001000010001","001000010001","000100010001","000100010001","000100010000","000100010001","001000010001","000100010001","000100010000","000100010001","000100010001","000100010000","001100100010","001000100001","000100010000","001000010001","010101000101","011001010110","010101000101","010000110011","001000100001","001000100001","011001010110","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000100010","001000100001","000100010001","000100010000","010000110011","010101010101","010101000100","010000110011","001000100010","001000100001","010101000101","011101100111","011101100111","011101100111","011101100111"))
	-- 4
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001001","100001111001","100001111001","100110001010","101010011011","101010011011","101010011100","101010101100","101010011100","101010011100","101010011011","100110011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001010","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011100","101010011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100101111000","100101100111","100101100110","100001100110","100101110111","100101110111","100101111000","100110001001","100110001010","101010011011","101010101100","101010011011","100110011010","100010001001","100110001001","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100101110111","100001010100","011100110011","011000110010","011000100010","011100110011","011101000011","011101000100","100001111000","100110001001","100110001010","101010011011","100110001010","100110001001","100110001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100101111000","100001000100","011100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011001000101","100110001001","100010001010","100110001001","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100101110111","011000110011","010000100001","010000100010","010100100010","010100110011","011001000100","011000110100","010100100010","011000110011","100110001010","100110001010","100110001010","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100101111000","011101000011","010100110010","011000110011","011101000101","100001010110","100101100111","100101100110","011000110011","010100100010","100101111000","100110001010","100110001001","100110001010","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110001001","100001010101","011101000101","100001010101","100001010101","100001010110","100101100111","100101100111","011101000101","010100110011","100001100111","100010001001","100110001001","100110001001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110001010","100001010110","100001010101","100001010101","100001010101","100001010101","100001010110","100001010110","100001010110","011000110011","100001100111","100110001001","100110001001","100001111001","100001111000","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","100101100111","011101000101","011000110100","011101000100","100001010101","011101000100","100001010110","100101010111","011101000101","100001010110","100110001010","101010011010","100110001010","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","100110001001","011101010101","011000110011","011101000100","100101010110","100001010110","100001010111","100101010111","100101010110","100001010110","100110001010","100110011010","101010011010","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001001","100110001010","100001010110","011101000100","011101000100","100001010110","100001010110","100001010110","100101010111","100001010110","100101111000","101010011011","101010011010","101010011010","100110011010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110011010","100010001001","100010001001","100010001001","100001100110","011101000100","011101000100","100001010101","100001010110","100001010110","100001010110","100001010110","100101111000","100110001010","100110011010","100110001010","100110011010","100110011010","101010011010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100001111001","100101111001","011101000101","011101000100","011101000101","100001010110","100001010110","100001010110","011001010101","011001010101","100101111001","101010011010","101010011010","100110001010","100110001010","100110001010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100001111001","100001111000","100001111000","100110001010","101010011011","100001100111","011101000100","011101000100","100001010101","100001010110","100001010110","011001010101","011001010101","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001","100110001001","100110001010","101010011011","100110011010","100010001001","100001111000"),
		("100001111001","100001111000","100001111000","100001111000","100110001001","101010011011","101010011010","100001010101","011101000100","100001000101","100001010101","100001010110","011001000101","011001010101","011001010110","011001010101","011001010110","011001010110","011001010110","011001010110","011001010110","011101100110","011101101000","100110001010","101010011011","100110001010","100001111001"),
		("101010011011","100110001001","100001111000","100001111000","100001111001","100110001010","100110001010","100001010110","011000110011","011000110011","011101000100","100001010101","011001000101","011001010101","011101100111","001100100011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100011","011001010110","100110011010","100110001010","100001111001"),
		("101010011011","100110001001","100001111000","100001111000","100001111001","100001111001","100001100111","011101000101","011000110011","011000110011","011101000100","100001010101","011001010101","011001010110","100001111001","010001000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100001111001","100001111000"),
		("101010011010","100110001001","100001111000","100001111000","100001111001","011101100111","010000110011","011001000101","011101000101","011000110011","011101000100","100001000101","011101010110","100001110111","100110001001","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010101000100","100001111001","100001111001"),
		("101010011010","100110001001","100001111000","100001111000","011001010101","001100100010","001000100010","010001000100","100001111000","011101000101","011101000100","100001010101","100001100111","100001111000","100110001001","010101010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","010000110011","100001111001","100001111000"),
		("101010011010","100110001001","100001100111","010100110100","001100100010","001000100001","001000100001","001100100010","011101100111","100001111001","100001010111","100001010110","100001100111","100001111000","100110001001","010101000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100001111001"),
		("101010001010","011101010110","010000100010","001000100001","001000100010","001000100010","001000100010","001000100010","011001010110","100001111001","100001111001","011101100111","011101100110","011101100111","100001111000","010001000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","010000110100","100001111001"),
		("011001000101","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110100","011101100110","010101010101","010101000101","010101000101","011001010101","011001010110","010001000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","100001111000"),
		("001000100001","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","010101000100","011001010101","011001010101","011001010101","011001010110","010101000100","001100100010","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","010000110011"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","011001010101","011001010101","011001010101","011001010110","010101000100","001100100010","001000100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001"),
		("001000100001","001000100001","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","011001010101","010101010101","010101010101","011001010101","010101000100","001100110011","001000100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001100100010","010101000101","010101010101","011001010101","010101010101","010101000100","010000110011","001000100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000010001","001000100001","001000100001"),
		("001000100001","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","010001000100","010101000101","011001010101","010101010101","010101000100","010000110011","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000010001","001000100001","001000100001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100001","001000100010","001100110011","010101000101","011001010101","010101000101","010001000100","010000110011","001100100010","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000010001","001000010001","001000100001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001100100010","010101000100","011001010101","010101000100","010001000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000100010","001000100010","001000100010","010000110100","010101000101","010001000100","010000110100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000010001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001000100010","001100110011","010101000101","010001000100","010000110100","010000110100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","010000110100","001000100010"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001100110011","010101000100","010001000100","010000110100","010000110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001"),
		("001000100001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001100110011","010101000100","010000110100","010000110100","010000110011","010000110011","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000010001","001000100001","010000110011"),
		("001000010001","000100010001","000100010001","000100010000","000100010000","000100010001","000100010000","000100010001","001000010001","001000010001","001000100001","001000100001","001100110011","010000110011","010000110100","010000110011","010000110011","010000110011","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","011000110100","011000110011"),
		("001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","001000010001","000100010001","001000010001","001000100001","001100110011","001100110011","010000110011","010000110100","010000110011","010000110011","001100100010","001000100001","001000100010","001000100010","001000100001","001100100010","001100100010","011000110011","011000110011"),
		("001000010001","000100010000","000100010000","000100010000","000100010000","001000010001","001000100001","000100010001","001000010001","000100010000","001000010001","001000010001","001100110010","001100100011","010000110011","010001000100","010000110100","010000110011","001100100010","001000100001","001000100001","001000100010","001000100001","001000010001","001000010001","010100110011","011101000101"),
		("001000010001","000100010001","000100010001","000100010001","001100100010","001000100001","001000100010","001000100001","001000010001","000100010001","000100010000","001000010001","001100110011","001100100010","001100100011","010000110011","010000110011","010000110011","001100100010","001000100001","001000100001","001000100010","001000100001","000100010000","001000100001","011000110100","011101000101"),
		("001000010001","001000010001","001000010001","001000010001","011001000101","001100110010","000100010000","001000100001","001000010001","001000010001","000100010000","001000010001","001100110011","001100100010","001100100010","001100110011","001100100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","000100010000","001000010001","001100100010","010100110011"),
		("001000010001","000100010001","001000010001","000100010001","001000100010","001100100010","000100010000","000100010000","000100010001","001000010001","000100010000","000100010000","001100100010","001100100010","001000100010","001000100010","001100100010","001100100010","010000110011","010000110011","001100100010","001000100010","001000100001","000100010001","000100010001","001000100001","001000100010"),
		("001100100010","001000100001","001000010001","000100010000","001000010001","001000100001","000100010000","000100010000","001000010001","001000010001","000100010000","000100010000","001100100010","001100100010","001000100010","010001000100","010101000101","010101010101","011001010101","010101000101","010000110011","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010"),
		("001100100010","001000010001","000100010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","000100010000","000100010000","001100100010","001000100010","001000100010","010101010101","011001010110","011001010101","011001010101","010101010101","010000110100","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("001000100001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000100010","001000100001","001000010001","010001000100","011001010101","010101000101","010101000101","010101000101","010000110100","001100100011","001000100001","001000100010","001000100010","001000100010","001000100010"))
	-- 5
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011100","101010101100","101010011100","101010011100","101010011100","101010011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001001","100110001010","100110001001","100001111001","100110001001","101010011011","101010101100","101010101100","101010101100","101010011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","101010011010","100110001001","100110001001","100110011010","101010011011","101010101100","101010011011","100110011010","100110001001","100110001010","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011100","101010001001","100101110111","100001010101","100001010101","100001010110","100101110111","100110001010","101010011011","100110001010","100110001001","100110001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101010101100","100101111000","100001010100","011101000011","010100100010","010100100010","011000110010","011101000011","011101010101","100101111001","100110001001","100110011010","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101010011011","100001010100","011000110010","010100100010","010100100010","010000100010","010100100010","010100100010","010100100010","011101010110","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101010001010","011101000100","010100100010","010100100010","010100110010","011000110100","011101000100","011101000100","010100100010","011001000100","101010011010","101010011011","101010011010","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101010001001","100001010100","011101000100","011101000100","100001010101","100101100110","100101100111","100101100111","011000110100","010100110011","100101111001","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110011011","100101111000","100001000101","100001010101","100001010101","100001010110","100101010110","100101100111","100101100111","100001000101","011000110011","100001111000","100001111001","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110011011","100101111000","011101000101","100001000101","011101000100","100001010101","100001010110","100001010101","100001010110","100001010110","011001000100","100110001001","100001111001","100001111000","100001111001","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010101100","100110001010","100110001010","101010011011","101010011011","100110001010","100001100110","011101000100","011000110100","011101000100","100001010110","011101000101","100001010110","100101010110","011101000101","100110001001","100110001001","100001111001","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100101111000","100001010101","011101000100","011101000101","100101010111","100001010110","100101010111","100101010111","100001010110","100101111000","101010011010","100110001010","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110011010","100010001001","100110001001","100110001001","100110001010","101010011011","100101111000","100001010101","011101000100","011101000100","100001010110","100001010110","100101100111","100001100111","100001010111","100110001001","101010011010","100110011010","101010011010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100110001010","100110011010","101010101100","100110001001","100001010110","011101000100","011101000100","100001010101","100001010110","011001010101","011101010110","100101111000","101010011010","100110011010","100110001010","100110001010","100010001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100010001001","100010001001","100001111001","100001111001","100110001010","101010011011","101010101100","101010011010","100001100111","011101000100","011100110011","011101000100","011101010101","011001010101","011101010110","100110001001","101010011010","100110001010","100001111000","100001111000","100001111000","100010001001","100110001010","101010011011","100110011010","100010001001","100001111000"),
		("100010001001","100001111000","100001111001","100001111000","100110001010","101010011011","101010011011","100110001010","100001111000","100001010110","011101000100","011101000101","011101010101","010101000101","011101010110","100101111001","100110001010","100110001001","100001111000","100001111001","100110001001","100001111000","100001111001","100110001010","101010011011","100110001010","100001111001"),
		("101010011011","100110001001","100001111001","100001111001","100001111001","100110011010","100110001010","100001111000","100001111001","100001110111","011101000100","011101000100","011001010101","010101000101","011101010110","100101100111","100001111000","100001111000","100001111001","100110001010","101010011010","100110001001","100001111000","100010001001","100110011010","100110001010","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100010001001","100001111001","100001111001","100001111000","100110001001","100101111000","011100110100","011100110011","011101010101","011001010101","011101010110","100001010111","011101010110","010000110011","011001010101","011101100111","100001111000","100110001001","100001111000","100001111001","100110001010","100001111001","100001111000"),
		("101010011011","100110001010","100001111001","100001111000","100001111001","100001111000","100001111000","100110001001","100110001010","100101111000","011101000100","011100110100","011101000101","011101100111","100001100110","100001010110","100001111000","001100110011","001100100010","001100100010","001100100010","010000110011","010101000100","010101000101","011101100110","100001111000","100001111001"),
		("101010011011","100110001010","100001111000","100001111001","100110001001","100110001010","100001111001","100110001001","100001111000","100001100111","011101000100","011101000100","011101000101","100001111000","011101010110","100001100111","100010001001","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001100100010","001100110011","011001010110"),
		("101010011010","100110001001","100001111001","100010001001","100110001010","101010011010","100101111000","011001000101","010100110011","100001100111","100001100111","011101000100","100001010110","100001111000","011101010110","100001111001","100001111001","001100110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100110011"),
		("101010011011","100110001001","100010001001","100110001001","100110001001","100001100111","010100110011","001100100010","001100100010","011101100111","100010001001","100001100111","011101010101","011101100111","100001111000","100110001010","011101100111","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","100110001010","100110001001","100001111000","011101000101","010000100010","001000100010","001000100010","001000100010","011101010110","100001111000","100001111001","011101100110","011001010101","100001111000","100110001010","011001010101","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010"),
		("101010011011","100110001001","011101010110","010100110011","001100100010","001000100010","001000100010","001000100010","001000100010","010000110100","010101000101","010101000101","010101000101","010101010101","011001010101","011101100111","010101000100","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100101111000","010000110011","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","010101010101","010101010101","010101010101","011001010101","010001000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100001111000","001100100010","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101010101","010101010101","011001010101","011001010101","010101000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001"),
		("100110001001","100001111000","001100100010","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","010101010101","010101000101","010101000101","010101000101","010101000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001001","011101100111","001100100010","001000010001","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","001100110011","010101000101","010101000101","010101000101","010101000100","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001010","011101100111","001000100010","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100001","001000100010","001100100010","010101000100","010101000101","010101000100","010101000100","010001000100","001100100010","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001"),
		("100110001010","011001010110","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001000100010","010000110100","010101000101","010101000100","010000110100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001"),
		("100110001001","011001010110","001000100001","001000010001","001000010001","001000010001","001000010001","000100010000","001000100001","001000100010","001000100010","001000100001","010000110011","010101000101","010101000100","010001000100","010001000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000010001"),
		("100110001001","011001010110","001100100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001000100010","001100100010","010101000100","010101000100","010000110100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001100110011","001000100010"),
		("100110001001","011101100110","001100100010","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001100100010","010101000100","010101000100","010001000100","010000110100","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001"),
		("100110001001","011101100110","001100100010","001000010001","000100010001","001000010001","000100010001","000100010000","001000010001","001000100010","001000100001","001000100010","001100100010","010101000100","010101000100","010001000100","010000110100","001100110011","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000010001"),
		("100110001001","011101010110","001000100010","001000100001","000100010000","000100010001","000100010001","001100100001","010000110010","010100110011","010000110011","001000100010","001100100010","010000110100","010001000100","010001000100","010000110011","001100110011","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001"),
		("100110001001","011101010110","001000100001","001000010001","000100010000","000100010000","001100100010","011101010101","100001010101","100001010101","011000110100","001000100010","001000100010","010000110100","010000110100","010001000100","010000110011","010000110011","001000100010","001000100001","001000100010","001000100010","001000100001","001000100010","001000100001","001000100001","000100010001"),
		("100110001001","011001010110","001000100001","001000010001","000100010001","001000100001","010100110011","011101000100","011000110011","011101000100","100001000101","001100100010","001000100010","010000110100","010000110100","010000110011","010000110011","010000110011","001100100010","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","000100010001"),
		("100110001001","011001010110","001100100010","001100100010","001000100010","001100100010","010000100010","011000110100","011000110011","011101000100","100001010101","001100100010","001000100010","010000110011","010000110011","010000110011","010000110011","010000110011","001100100010","001000100001","001000100001","001000100010","001000100010","001000100010","001100100010","001100100010","001100100010"),
		("100110001001","011101100111","001100100011","001000100010","001100100010","001000100010","001000100001","010100110011","011100110011","011101000100","011101000100","001100100010","001100100010","010000110011","010000110011","010000110100","010000110011","010000110011","001100100010","001000100001","001000100001","001000100010","001000100001","001100100010","011001000100","011101000100","100001000101"),
		("100001111000","100001111000","010101000100","001000100010","001000100010","001000100010","001000100010","010000100010","011000110011","011000110011","010000100010","001000010001","001100100010","010000110011","001100110011","010000110011","010000110011","010000110011","001100100010","001000100001","001000100001","001000100001","001000010001","010000100010","011000110100","011101000101","100001010110"),
		("100001111000","100001111000","011101100110","001100100010","001000100010","001100100010","001100100010","001000010001","001000100001","001000010001","000100010000","000100010000","001100100010","001100110011","001100100010","010000110011","010000110011","001100100010","001000100010","001000100001","001000010001","001000010001","000100010001","001100100010","011000110011","011101000100","100001010101"),
		("100001110111","100001110111","011101100111","010101000100","010001000100","010000110011","001100100010","001000100001","001000010001","001000010001","000100010000","000100010000","001000100001","001100110011","001100100010","001000100010","001000100001","001000100010","001100100010","001100100010","001000010001","000100010000","001000010001","000100010000","001100100010","010100110011","011101000100"),
		("011001100110","011001010110","011101100110","011101100110","011101100111","011101100110","011001010101","010101000100","001000010001","000100010000","000100010000","000100010000","001000010001","001100100010","001000100010","001000100001","001100100010","001100110011","001100110011","001100110011","001000100001","000100010001","001000010001","000100010000","000100010000","001100100010","010100110011"))
	-- 6
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001100111","100001111000","100001111000","100001111001","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","101010011010","100110001010","100110001010","100010001010","100010001010","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111000","100001111001","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011100","101010011100","101010011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110011010","101010011011","101010101100","101010101100","101010011100","101010101100","101010011100","101010011011","100110011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100001111001","100001111001","100110001001","101010001001","101010001000","100110001000","101010001010","101010011011","101010101100","101010011100","101010011011","100110001010","100110011011","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001001","100110001010","100101111000","100101010101","100001010100","011000110011","011000110010","011000110011","100001010101","100101111000","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","100001010101","011100110011","011000110010","010100100010","010100100010","010100100010","011000110010","011000110011","100001100111","100110001010","100110011011","100110001011","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010101100","101010101100","101010011010","100001010101","010100100010","010000100001","010100100010","010100100010","010100110010","010100110011","010100100010","011101010101","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101110101100","101110101100","101110101100","101010001001","100001000100","011000110011","011000110011","011101000100","100001010101","100001010110","100001010110","011000110011","011001000100","101010011011","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101100","101110101101","101110101101","100110001001","100001000100","100001010101","100001010101","100001010110","100101100110","100101100110","100101100111","100001000101","011000110100","100110001010","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","100101111000","011101000100","100001010101","100001010101","100001010101","100001010110","100101010110","100101010111","100001010110","011001000100","100110011010","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011010","100001010101","011101000100","011100110100","011101000101","100001010101","011101000101","100001010110","100001010110","011101010101","100110011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110001011","101010011011","101110101100","101110101100","101010011011","100101111000","011101000101","011101000100","011101000100","100001010110","100001010110","100001010110","100101010111","100001010110","100110001001","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110001010","100110011011","101010101100","101110101100","101010011010","100101100111","100001010101","011101000100","011101000101","100001010110","100101100110","100101100111","100101010111","100001010111","100001111001","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001011","100110001010","100101100111","100001010110","011101000100","011101000100","100001010110","100101010111","100101010111","100101010111","100001101000","100001111001","100110001001","101010011011","100110011011","100010001001","100001111001","100110001010","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110011011","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100101110111","011101000100","011101000100","100001010101","100001010110","100101010110","100101100111","100110001001","100110001010","100110001001","100010001010","100001111001","100001111001","100001111001","100110001010","100001111001"),
		("101010011011","100110011011","100010001001","100110001001","100110001010","100110001010","101010011011","101010101100","101010011011","100110001010","100110001010","100110001001","100001010110","100001010110","100001010110","100001010111","100101010111","100101100110","100101111001","101010011010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","100110001010","100001111001","100001111001","100110001010","100110011010","101010101100","101010101100","101010011011","100110001001","100001111001","100110001001","100001111000","011001010101","011101010110","100001100110","100001010110","100001010110","100101101000","011101100111","100001111001","101010011011","101010011011","101010011011","100110001010","100001111001","100001111000"),
		("100010001001","100110001001","100001111001","100001111001","100110001010","101010011011","101010101100","101010011011","100101111001","100001111000","100001111000","100001111000","011101100111","011001010101","011101010110","100001010101","100001010110","100001010110","100001100111","010101000100","010000110011","011001010110","100001111000","100110001001","100110001010","100010001001","100001111001"),
		("100110001001","100001111001","100001111001","100001111000","100110001010","101010011011","101010011011","100110001010","100001111000","100110001001","100110001010","100001111001","100001100111","011001000101","011101010110","100001010101","100001010110","100001010110","100001111000","010101000100","001100100010","001100100010","001100100010","010000110011","010101000100","011001010110","011101100111"),
		("101010011011","100110001010","100001111001","100001111001","100010001001","100110011010","100110001010","100001111000","100001111001","100110001010","100110001010","100110001001","011101100110","010101000101","011001010101","011101010101","100001000101","100001010110","100110001001","010101000100","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010"),
		("101010011011","100110001010","100001111001","100010001001","100010001001","100001111001","100001111001","100001111000","100010001001","100110001010","100101111001","011101100110","100001100111","011001010110","011001010101","011101000101","011101000101","100001111000","100001111001","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","100001100111","010100110011","010100110011","100001111000","100001111000","011101010101","011101000100","100001100111","100110001010","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111000","100001111001","100110001001","100110001010","100001111001","100110001001","011101010110","010000110011","001100100010","001100100010","100001100111","100001111000","011101100111","011101010110","100001100111","011101111000","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001001","100001111001","100010001001","100110001010","101010011010","100101111000","011001000101","010000100010","001000100010","001000100010","001000100010","011001010101","100001111000","011001010110","011001010101","011001010101","010101000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100110001001","100110001010","100101111000","010100110011","001100100010","001100100010","001000100010","001000100010","001000100001","001100100010","011101100110","011001010110","010101010101","010101010101","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100110001001","100110001001","011101100111","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","010001000100","010101000101","011001010101","010101000101","001100110011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010"),
		("101010011011","100110001001","100010001001","100110001001","100110001001","011101100110","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101000101","010101010101","010101000100","001100100011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100110001001","101010011010","011101100111","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010001000100","010101000101","010101000101","010101000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","101010011010","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","010001000100","010101000100","010101000101","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001"),
		("100110001001","100010001001","100110001001","100110001001","100110001001","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110100","010001000100","010101000101","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100010001001","100010001001","100010001001","100110001001","100001111001","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","010000110011","010101000100","010000110100","010000110011","010100110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001001","100110001001","100110001001","100110001001","100110001010","100001111001","001100100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","010000110011","001100110011","010000110100","010000110011","010100110100","100001000101","011101000100","010100110011","001100100010","001000100010","001000100010","001000100001","001000010001","001000100001"),
		("100110001010","100010001001","100110001001","100110001001","100110001010","100110001001","010000110010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","001100100010","010000110011","010000110011","011101000101","100001010101","100001010101","100001010101","010100110011","001000100010","001000100010","001000100001","001000010001","001000010001"),
		("100110001001","100110001001","100010001001","100110001001","100110001010","100110001010","010000110011","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","010000110011","001100100010","010000110011","010000110011","011001000100","011101000100","100001010101","100001010101","100001000101","010000100010","001000100001","001000100001","001000100001","001000010001"),
		("100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","010101000100","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","010000110011","001100100010","010000110011","010000110011","010100110011","011101000100","100001000101","100001010101","100001010101","011001000100","001000100001","001000100010","001100110011","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","100110001001","100101111001","010101000100","001000100001","001000010001","001000100001","001000100001","001000100010","001000100001","010000110011","001100100010","010000110011","010000110011","010000110011","011000110011","100001000101","100001010101","100001010101","011001000100","001000100010","001000100010","001100100010","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","100110001001","100101111000","011001000101","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","001100100010","010000110011","010000110011","001100100010","010000100010","011000110011","011101000100","100001000101","011001000100","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100110001001","100101111000","100101111000","100001100111","010101000100","001100100010","001000100001","001000010001","001000010001","001000100001","001000100001","010000110011","001000100010","001100110011","001100100010","001000100010","001000100001","001000100001","001100100001","010000100010","001100100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100101111001","100001100111","100001000101","011101000100","010100110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","010000110011","001000100010","001100100010","001100100011","001100100010","001000100010","001000100001","001000010001","000100010000","001000010001","001000100010","001100100010","001000100010","001000100010"),
		("100110001001","100001110111","100001010101","100001010110","011101000101","010100110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","001000100001","001000100010","001100100010","001100100010","001000100001","001000100001","001000010001","000100010000","001000010001","001100100010","001100100010","001000100001","001000100001"),
		("100110001001","100001111000","011101000101","100001010110","100001010101","011000110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000010001","000100010000","000100010001","001000010001","001000010001","001000010001","001000010001"),
		("100010001001","100001111000","011101010110","011101000101","100001000101","011000110011","001000100001","000100010001","000100010000","000100010001","001000010001","001000010001","001000100001","001100110011","001100100010","010000110100","010001000100","010001000100","010000110011","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100010"),
		("100001111000","100001111000","011101010110","011000110011","011000110011","001100100010","001000100001","001100110011","010101000101","001100110011","000100010000","001000010001","001000010001","001100110011","001100100010","010101000100","010101010101","010101010101","010101000100","001000100001","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","011101100110","010000110011","010000110011","010101000101","011101100110","100001111000","100001111000","010001000100","001000010001","000100010000","001000010001","001100110011","001100100010","010101000101","010101000101","010101010101","010101000100","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100001110111","100001110111","100001100111","011101100111","100001111000","100001111000","100001111000","100001111000","011001010110","010101000100","001000010001","000100010000","001000010001","001100100010","001100100010","010101000101","010101000101","010101000101","010101000100","001100100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("011001100110","011001100110","011101100110","011101100110","011101100111","011101100110","011101100111","011001010110","010000110011","001000100001","000100010000","000100010000","001000010001","001100100010","001100100010","010101000100","010101000100","010101000100","010101000100","001100100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"))
	-- 7
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100010001001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100101100110","100001010101","100001010100","011101000011","011101000100","100001100111","100110001001","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111001","100001100111","011100110011","011000110010","010100100010","010100100010","010100100010","011000110010","011101000100","100101111001","100010001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100101111001","100101010101","011000110010","010000100001","010000100001","010100100010","010000100001","010100100010","010100100010","011101000101","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100101111000","100001010100","011000110011","011000110011","011000110011","011000110011","011001000100","011000110100","010100100010","011000110011","101010011010","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100001111001","100001111001","100101100110","100001000100","100001000101","100001010101","100001010110","100101100110","100101100111","100101100111","011001000100","011000110100","100110001010","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001001","100110001010","100110001001","100001010101","011101000100","100001010101","100001010101","100001010110","100101100110","100101100111","100101100111","011101000101","011000110100","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","101010011011","100101100111","100001000101","011101000100","011101000100","100001010101","100001010101","100001010101","100001010110","011101000101","011101000101","100110001010","100010001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010101100","101010101100","101010101100","101010011100","100110001001","100001100110","011101000100","011101000100","011101000101","100001010110","011101000101","100001010110","100001010101","100001100111","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101110101100","101110101100","101110101100","101010011100","101010011011","100101100111","100101100111","011101000101","011101000100","011101000101","100101010110","100101100110","100101100111","100001010110","100001100111","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101100","101110101101","101110101100","101010011011","101010011011","100101101000","100001100110","011101000101","011101000100","011101000101","100001010110","100101100111","100101010111","100101010110","100101111000","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","101010011011","100110001010","100101111000","100001010101","011101000100","100001000101","100101010110","100101010111","100101010111","100101101000","100110011010","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","101010011011","101010011011","100110001001","100001010101","011101000100","011101000100","100001010110","100001010110","100101010110","100110001010","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110001011","101010011011","101110101100","101110101100","101010101100","101010011011","100110001010","100001111001","100001100110","100001000101","100001010101","100101100110","100101010111","100001010110","100110001001","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110001010","100110011011","101010101100","101110101100","101010011011","100110001010","100001111001","100001111001","100001100110","011101000100","011101000100","100001000101","100101010110","100101010111","011101100110","011101100111","101010011010","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100001111001","100110001001","100001100111","011101000100","011101000100","100001010110","100101010111","100101100111","011001010110","001100100010","011001010101","100001111000","100001111000","100001111001","100110001010","100010001001"),
		("101010101100","101010011011","100110001010","100110001010","100110011011","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100110001010","100110001010","100001010101","011101000100","011101000100","100001000101","100001010110","100101111001","011001010110","001100100010","001100100010","010000110011","010000110011","011001000100","011001010101","011001010110"),
		("101010011011","100110011011","100010001001","100110001001","100110001001","100110001010","101010011011","101010101100","101010011011","100110001010","100110001001","100110001001","100101111001","100001010110","100001010110","100001010101","011101000100","100001100111","100110001010","010101000101","001100100010","001000100010","001000100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100110001010","100110001010","100110011010","101010101100","101010101100","101010011011","100110001001","011101100110","011101010101","100101111000","100001100111","011001010101","011101010101","100001010110","100110001001","100001111000","001100110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010101100","101010011010","100001111000","011001000100","010000100010","010100110011","100101111000","011101100111","011001000101","011101100110","100001111001","100110001010","010101000101","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100001111001","100001111001","100001111000","100110001010","101010011011","101010011010","100001100111","010100110011","001100100010","001100100010","010000110010","100001100111","011101010110","011001010101","011001010110","011001010110","011001010101","001100100011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111001","100010001001","100110001010","011001010101","010000100010","001100100010","001000100010","001000100010","001000100010","010000110011","011001010101","011001010101","011001010110","011001010101","010001000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100010001001","100110001001","100001111000","010000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","011001010101","011001010101","010101010101","010000110011","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100010001001","100001111001","100001111001","100001111000","010000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","011101100111","011001010101","010101000101","001100110011","001000100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111001","100110001001","100001111000","010000100010","001000100010","001000100001","001000100010","001100100010","001100100010","001000100010","010101000101","100001100111","011001010101","010101000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001001","100001111001","100010001001","100110001010","100110001001","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000101","100001111000","010101000101","010001000100","001100100010","001100100010","001100100011","001100100010","001100100010","001100100010","001000100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100110001001","100110001010","100110001010","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","011001010110","010101000100","010000110011","011001000100","100001010101","100001010101","011101000101","010100110011","001000100010","001000100010","001000100010","001100100010","001000100010"),
		("101010011011","100110001010","100010001001","100110001001","100110001001","100110001010","010100110100","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","010000110011","010101000101","010001000100","001100100010","011001000100","100001000101","100001000101","100001000101","100001000101","010000110011","001000100010","001000100010","001100100010","001000100010"),
		("101010011011","100110001001","100010001001","100110001001","100110001001","100101111001","010100110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101000101","010000110100","001100100010","010000110011","011101000101","100001000101","100001000101","100001010110","100001000101","001100100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100110001001","101010011010","100101111001","010101000100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101000100","010000110011","001100100010","001100100010","011100110100","011101000100","100001000101","100001010110","100001010110","010000110011","001000100001","001000100010","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","100110011010","100101111000","011001000101","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","010000110100","010101000100","010000110011","001000100010","001000100010","001100100010","010000100010","010100110011","011101000101","100001010110","010100110011","001000100001","001000100001","001000100001"),
		("100110001001","100010001001","100110001001","100110001001","100001111001","100101111000","100001100111","001100100011","001000100010","001000100010","001000100010","001000100010","001000100010","010000110100","010101000100","010000110011","001000100001","001000100001","000100010001","000100010000","000100010000","010000100010","010100110011","010000100010","001000100010","001000100001","001000100001"),
		("100110001001","100110001010","100010001001","100110001001","100001111000","100110001001","100110001001","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011","010101000100","001100110011","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010001","000100010001","001000100001","010000110011","010001000100"),
		("100110001010","100110001010","100110001001","100110001001","100110001001","101010011011","100110001010","010001000100","001000100001","001000100001","001100110011","001000100010","001000100001","010000110011","010101000100","001100100010","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001000010001","001100100010","001100110010"),
		("100110001010","100110001001","100110001001","100110001001","100110001001","101010011010","100101111001","010000110011","001000100010","001100100010","010000110100","001000100010","001000100010","010000110011","010101000100","001100100010","001000100001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001"),
		("100110001001","100110001001","100010001001","100110001001","100110001010","101010011010","011101100111","001100100010","001000100001","001100100010","010000110011","001000100010","001000100010","010000110011","010000110011","001000100010","001000010001","001000010001","001000010001","001000010001","000100010000","001000100001","001100100010","001000010001","001000010001","001000010001","001000010001"),
		("100110001001","100110001001","100110001001","100110001001","100001100111","100001010110","010100110011","001000100001","001000100001","001000100001","001100100010","001000100001","001000100001","001100100011","010000110011","001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000100001","001000010001","000100010001","001100110010","001000100001"),
		("100110001001","100110001001","100010001001","100001100111","100001000101","011101000100","010100110011","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001100110011","010000110011","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010"),
		("100110001001","100110001001","100001111000","100001010110","100001010110","100001010101","011000110011","001000100001","001000010001","001000010001","001000100001","001000010001","001000010001","010000110011","001100110011","001000010001","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100110001001","100101111000","100001010110","100001010110","100001010110","011000110100","001000010001","001000010001","001000100010","001000100001","001000100001","001100100010","010101000100","010000110011","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001001","100110001001","100001100111","100001000101","100001000101","011000110011","010001000100","011101100111","011001010101","001000010001","001000010001","001100100010","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100010001001","100001111000","011101000101","011101000101","011101100111","100001111001","100110001001","010001000100","000100010001","001000010001","001100110010","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001001","100010001001","100010001001","100010001001","100110001001","100001111001","100001111000","100001111000","100001111000","001100100010","000100010001","001000010001","001100110011","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100010001001","100001111001","100001111000","100001111001","100110001001","100001111000","100001111000","100001111001","011101100111","001000100010","000100010001","001000010001","010000110011","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100110001001","100110001001","011001010110","001000100001","001000010001","001000010001","010000110011","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","100001110111","100001111000","100001111000","100001111000","100001111001","100001111001","010000110100","001000100001","001000010001","001000010001","010000110100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100001110111","100001100111","100001100111","100001100111","100001111000","100001111000","100001111000","011101100111","010000110011","001000100001","001000010001","001000010001","010100110100","010101000100","010000110011","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100001","001000100010","001000100010"),
		("011001100110","011001100110","011101100110","011101100110","011101100111","011101100110","011101100111","010101010101","001100100010","001000010001","000100010000","001000100001","010000110100","010000110011","010000110011","001000100010","001000100001","001000010001","001000100001","001000100001","001000100001","001000100010","001000100001","001000100010","001000100001","001000100010","001000100010"))
	-- 8
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100010001001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100001111000","100101010101","100001010100","011101000100","011101000100","011101010101","100001111000","100110001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111001","100001111000","100101100110","011000110010","010100100010","010100100010","010100100010","010100100010","011000110011","100001100111","100010001010","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100001111001","100101100111","100001000100","010100100010","010000100001","010000100010","010000100001","010000100010","010100100010","011000110011","100101111000","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100110001001","100101100110","100001000100","011000110011","011000110011","011000110011","011000110011","011000110011","010100110010","010100100010","100001111000","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100001111001","100001111001","100101111000","011101000100","100001010101","100001010101","100001010110","100101010110","100101100111","100101100110","100001010101","010100100010","100001111000","100110011011","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001001","100110001010","100110001001","100001100111","011101000100","100001010101","100001010101","100001010110","100101100110","100101100111","100101100111","100001010110","011000110011","100001100111","100010001010","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","101010011011","100101111000","100001010101","100001010101","011100110100","011101000100","100001010101","100001010110","100001010110","100001010110","011000110100","100001111001","100110001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010101100","101010101100","101010101100","101010011011","100101111000","100101100111","011101000101","011101000100","011101000100","100001010110","011101000101","011101000101","100001010101","011101010110","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101110101100","101110101100","101110101100","101010101100","101010011011","100001010110","100101100110","100001000101","011101000100","011101000100","100001010110","100101100110","100101100110","100001010110","100001101000","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101100","101110101101","101110101100","101010011011","101010011011","100101111000","100101100110","011101000101","011101000100","011101000100","100001010110","100101010110","100101010111","100101010110","100101111000","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","101010011011","101010011010","100101111000","100001010101","011101000100","100001000101","100001010110","100101010111","100101010111","100101100111","100110001010","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","101010011011","101010011011","100110001001","100001010101","011101000100","011101000100","100001010110","100001010110","100101100111","100110001010","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110001011","101010011011","101110101100","101110101100","101010101100","101010011011","100110001010","100001111000","100001010101","011101000101","100001010101","100101010110","100101010110","100101100111","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110001010","100110011011","101010101100","101110101100","101010011011","100110001010","100001111001","100001100111","011101000100","011101000100","011101000100","100001010101","100101010110","100101100111","100001111001","100110001010","101010011010","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100001111001","100001100110","100001000101","011101000100","100001010101","100001010110","100101010111","100001100111","011001010101","100110001001","101010011010","100110001010","100001111001","100001111001","100110001001","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110011011","100110001010","100110001010","100110001010","100110001001","100001111001","100010001001","100101111000","100001000101","011101000100","011101000100","100001000101","100001010101","100101100111","011101100110","001100100010","010001000100","011101100110","100001100111","100001111000","100001111001","100110001001","100001111001"),
		("101010011011","100110011011","100010001001","100110001001","100110001010","100110001010","101010011011","101010011011","100001111000","011101010110","100001100111","100101111000","100001010110","100001010110","011101000101","011101000101","100001010110","100110001001","011001010110","001100100010","001100100010","001100100010","010000110011","010101000100","011001010101","100001100111","100001111000"),
		("101010011011","100110001010","100010001001","100110001010","100110001010","100110001010","100101111000","011101010101","010100110011","010100100010","100001010110","100101111000","011001010101","011001010101","011101010101","100001100110","100110001001","100010001001","010000110100","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","010000110011"),
		("100110001010","100110001010","100001111001","100010001001","100001100111","011001000101","010100110011","001100100010","001100100010","001100100010","100001010110","100101111000","011001010101","011001010101","100001110111","100110001010","100110001010","011001010110","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100001111001","100001111001","100001111001","010101000100","001100100010","001100100010","001000100010","001100100010","001100100010","010000110011","010101000100","011001010101","011001010101","011101010110","011101100111","100001111000","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111000","010000110011","001100100010","001000100010","001100100010","001100100010","001000100010","001000100001","010000110011","011001010101","011001010101","011001010101","011001010101","010101000101","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","100110001010","100010001001","100001111000","010000110011","001000100010","001100100010","001100100010","001000100010","001000100010","001000100001","010000110011","011001010101","011001010101","011001010101","011001010101","010001000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111000","010000110011","001000100001","001100100010","001000100010","001000100010","001000100010","001000100001","010000110011","011001010110","011101100110","011001010101","010101000101","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100001111001","100001111000","010000110011","001000100001","001100100010","001000100010","001000100001","001000100010","001100100010","010000110011","011101100110","011101100111","010101010101","010101000100","001100100011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001001","100001111001","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","011101100111","011101100111","010101000101","010101000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001100100010","001100100010","001100100010"),
		("101010011011","100110001010","100110001001","011101100110","001100100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100001","001100110011","011001010110","011001010101","010101000100","010000110100","001000100010","001000100010","001000100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001"),
		("101010011011","100110001010","100110001001","011101100110","001100100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100001","001100100010","010101000100","010101000100","010101000100","010000110011","001000100010","001000100010","001100100010","011101000100","011101000101","011001000100","010100110011","001100100010","001000100010","001000100010","001000010001"),
		("101010011011","100110001001","100001111001","011101100110","001100100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","010101000100","010001000100","001100100010","001000100010","001000100010","001100100010","011100110100","100001000100","100001010110","100001010110","011001000100","001000100010","001000100010","001000010001"),
		("100110001010","100110001001","100110001001","011101100111","001100100010","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010","010101000100","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","010100110011","011101000100","100001010110","100001010110","100001010101","010000110011","001000100001","001000100001"),
		("100110001001","100110001001","100110001001","011101100110","001100100010","001000100001","001000010001","001000100001","001000100010","001000100010","001000100001","001000100001","010000110100","010101000100","010000110011","001100100010","001000100001","001000100010","001000100001","001100100010","011100110100","100001000101","100001010110","100001010110","011001000100","001000100001","001000100001"),
		("100110001001","100010001001","100110001001","011101010110","001100100010","001000100001","001000100001","001000010001","001000100010","001000100010","001000100010","001000100010","010000110011","010101000100","010000110011","001000100010","001000100001","001000100001","001000010001","001000010001","010000100010","011000110100","011101000101","100001010101","011101000101","001100100010","001000100001"),
		("100110001001","100110001010","100110001001","011001010110","001100100010","001000100001","001000100001","001000010001","001000100001","001000100010","001100100010","001100100010","010000110011","010101000100","010000110011","001000100001","001000100001","001000100001","001000010001","000100010001","000100010001","000100010000","001100100001","011101000100","011101000100","001100100010","001000100010"),
		("100110001010","100110001010","100110001001","011101010110","010000110011","001100100010","001100100010","010101000100","011101010101","011101000100","011100110100","010100110011","010000110011","010101000100","001100110011","001000100001","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010000","001000010001","001000100001","001000010001","001000100001"),
		("100110001010","100110001001","100110001001","100001111000","010000110011","001100100010","010101000100","100001010110","011101000100","011100110011","011100110011","010100100010","010000110011","010101000100","001100110011","001000100001","001000100001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001"),
		("100110001001","100110001001","100110001001","100010001001","010100110011","010000100010","001100100010","010100110100","011101000100","011100110011","011100110011","010100100010","010000110011","010101000100","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","000100010001","001000010001","001000010001","001000010001","001000010001"),
		("100110001001","100110001001","100110001001","100110001001","011101010110","001100100010","001000100010","010000100010","011100110011","011000110011","011000110011","010000100010","010000110011","010001000100","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","001100110010","001000100001"),
		("100110001001","100110001001","100110001001","100110001001","100001111001","011101010110","010100110100","001100100001","010100110011","011000110011","010100100010","001000010001","010000110011","010000110100","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001"),
		("100110001001","100110001001","100110001001","100110001001","100110001010","100101111001","100001100111","010100110011","001100100001","001000100001","001000100001","001000010001","001100110011","010000110011","001000100010","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010"),
		("100110001001","100110001001","100110001001","100110001001","101010011010","100110001010","100101111000","100001111000","011001010110","001100110011","001000010001","001000010001","001100100010","001100100010","001000010001","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100110001001","101010011010","101010011010","100110001001","100001111000","011101100111","010000110011","001000010001","001000100010","010000110011","010000110011","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100010001001","100110001001","101010011010","101010011010","100001111001","100001111000","011101100111","001100110011","001000100001","010000110011","010101000100","010000110100","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100110001001","100010001001","100010001001","100010001001","101010011010","100110001001","100001111000","100001111000","011001010101","001100100010","001000100001","010000110100","010101000100","010101000100","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001"),
		("100010001001","100001111001","100001111000","100001111001","100110001001","100001111000","100001111000","100001111000","010101000100","001000100010","001000100010","010101000100","010101010101","010101000100","001000100010","001000100001","001000010001","001000010001","001000010001","001000100001","001100100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100110001001","011101100111","001100110011","001000100001","001000100010","010101000101","010101010101","010101000101","001100100010","001000100001","001000010001","001000010001","001000010001","001000100001","001100110011","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","100001110111","100001111000","100001111000","100001111000","100010001001","011001010110","001100100010","001000100001","001100100010","010101010101","010101010101","010101010101","001100110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001110111","100001100111","100001100111","100001100111","100001111000","100001111000","100001111000","011001010101","001100100010","001000100001","001000100010","010101010101","010101000101","011001010101","010001000100","001000100001","001000010001","001000010001","000100010000","000100010001","000100010001","001000010001","001000010001","001000100010","001000100001","001000100010","001000100010"),
		("011001100110","011001100110","011101100110","011101100110","011101100111","011101100110","011101100111","010101000100","001000100010","001000010001","001000100001","010101000101","010101000100","010101000101","010101000100","001000100001","001000010001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","001000100001","001000100010","001000100010"))
	-- 9
	,

		(	("100001111001","100001111001","100010001010","100001111001","100001111001","100010001010","100110001010","100110001010","100001111001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111001","100001111001","100010001010","100001111001","100110001010","100110001011","100110001010","100001111001","100001111000","100001111000"),
		("100010001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001001","100110001010","100110011010","100110001010","100110001001","100010001001","100010001001","100010001010","100010001010","100110001010","100110001010","100010001010","100001111001","100001111000"),
		("101010011011","100110011011","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001111001","100001110111","100101100110","100101100110","100001100110","100101110111","100110001001","100110001001","100110001001","100110001010","100010001001","100010001001","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100001111001","100101111000","011101000011","011000110010","011000110010","010100100010","010100100010","011000110011","100001100111","100110001001","100101111001","100110001001","100110001010","100110001010","100010001010","100001111001","100001111001"),
		("101010101100","101010011011","100110001010","100110011011","100110011011","100110011011","101010011011","101010011011","101010011011","100110001010","100001111001","100101100101","011000110010","010000100001","010000100001","010100100010","010100100010","010100100010","011100110011","100101111000","100110001001","100110011010","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("100110001010","100110011011","100110011011","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010","100010001001","100101110111","100001010100","011000110010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","100001010110","100110001001","100110001010","100110011010","100110001010","100010001001","100001111001","100001111001"),
		("100110001010","101010011100","101010011011","100110001010","100110001010","101010011011","100110001010","100010001010","100010001010","100110001010","100001100110","011101000011","100001000100","100001010101","100001010101","100001010101","100001010110","100001010101","010100110011","011101010101","100010001001","100001111001","100001111001","100001111001","100010001001","100110001010","100001111001"),
		("101010011011","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","011101000101","011101000011","100001010101","100001010101","100101100110","100101100110","100101100110","100101100111","011101000100","011101010110","100110001010","100110001010","100010001010","100001111001","100010001001","100110001010","100001111001"),
		("101010101100","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010101100","101010101100","101010011011","100001010110","011101000100","011101000100","011101000100","100001010101","100101010110","100101010110","100101100111","011101000100","100001100110","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010101100","101110111101","101010011011","100110011011","100110011011","101010011100","101110101100","101110101100","101110101100","101010011011","100101100111","100001000101","011101000100","011101000100","011101000101","100001010101","011101000101","100001010110","011101000101","100101111001","101010011011","101010011011","101010011011","100110011011","100010001010","100001111001","100001111001"),
		("100110011011","101010101100","101010011011","100110011011","100110011011","101010011011","101110101100","101110101101","101110101100","100101111000","100001010110","100101100110","100001000101","011101000101","100001000101","100101010110","100001010110","100101010110","100001100110","101010011010","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001"),
		("101010011011","100110011011","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","100110001001","100001010101","100001010110","100001000101","011101000101","011101000100","100001010110","100101100111","100101010110","100001100111","100110001010","101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101010011100","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101110101100","101010011011","100101111001","100001010110","011101000100","011101000100","100001010101","100101010110","100101010110","100001010110","100101111000","101010011011","101010011011","101010011011","101010011011","101010011011","100110001011","100001111001","100001111001"),
		("101110101101","101010101100","100110011011","100110011011","100110011011","100110001011","101010011011","101110101100","101110101100","101010101100","101010011011","100001010110","011101000100","011101000100","011101000101","100001010110","100101010110","100101100111","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001"),
		("101110101101","101010101100","100110001010","100110001010","101010011011","100110001010","100110011011","101010101100","101010101100","101010011011","100110001010","100001010110","011101000101","011101000101","100001010101","100101100110","100001010110","100001111000","100001111000","100001111000","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101100","101010011100","100110001010","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","100001111000","100001000101","011101000100","011101000100","100001000101","100001010110","100001010110","100101111000","100001111000","100001111000","100110001001","100110001010","100110001010","100001111001","100001111001","100110001001","100001111001"),
		("101010101100","101010011011","100110001010","100110001010","100110011011","100110001010","100110001010","100110001010","100010001001","100001111001","100001111000","100001000101","011101000100","011101000100","100001010101","100001010110","100001010110","100001111000","100110001001","100110001001","100001111001","100001111000","100001111000","100001111000","100001111001","100110001001","100001111001"),
		("101010011011","100110011011","100010001001","100110001001","100110001001","100110001010","101010011011","101010011011","100110001001","100101111000","100001100110","011101000101","100001010110","100001100110","100001010110","100001010110","100101100111","011001010101","011001010110","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000","100001111000"),
		("101010011011","100110001010","100010001001","100110001010","100110001010","100110001001","100101111000","011101010110","011101000101","100001100111","100001100110","011101000100","011001010101","011001010101","011101010101","100001010110","100101111001","010101000101","001100100010","010000110100","011001010110","100101111000","100110001010","100110001010","100110001001","100001111000","100001111000"),
		("100110001010","100110001010","100001111001","100001111000","100001100111","011001000101","010100110011","001100100010","001100100010","100001100111","100101111000","011101010101","011001010101","011001010101","011101100110","100001111000","100110001010","010101000100","001100100010","001100100010","001100100010","001100110011","010101000101","100001100111","100110001001","100010001001","100001111000"),
		("100110001010","100001111001","011101100110","011001000100","010000110011","001100100010","001100100010","001000100010","001100100010","100001100111","100110001001","100001111000","010101010101","011001000101","100001111000","100110001010","011101100111","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001100100010","010101000100","100001110111","100001111001"),
		("101010011011","100001111001","010000110011","001100100010","001100100010","001100100010","001000100010","001100100010","001100100010","011101010110","011101100111","011101100111","010101010101","010101010101","100001111000","100001111001","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","011101100111"),
		("101010011011","100001111000","001100100010","001000100010","001100100010","001000100010","001100100010","001100100010","001000100010","001000100010","010001000100","011001000101","011001010101","011001010101","011101100111","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100"),
		("101010011011","011101100111","001100100010","001000100010","001100100010","001000100010","001100100010","001000100010","001000100010","001000100010","010001000100","010101000101","011101010110","011101100110","011001010110","010001000100","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","010000110011"),
		("101010011011","011101100110","001100100010","001000100010","001100100010","001000100010","001100100010","001000100010","001000100001","001000100010","010101000100","010101000101","011101100110","011101100111","011001010101","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100011"),
		("101010011011","011001010101","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010001000100","010101000101","011101100111","011101100111","010101000101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001100100010","001100100010","001100100010"),
		("101010011011","010101000100","001000100001","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","010000110100","010101000101","011001010101","011001010110","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001100100010"),
		("101010011011","010101000100","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","010000110011","011001010101","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","010001000100","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","010000110011","010101000101","010101000100","010101000101","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","010000110100","001000100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100010","001000100010","001100110011","010101000101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100001","001100100010","010000110011","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","010000110011","001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001000100010","001000100010","001100100010","010101000100","010101000100","010001000100","001000100010","001000100010","001000100010","001000100010","001000100001","010000100010","011101000100","011000110011","010000100011","001000100010","001000100010","001000100001","001000100001"),
		("100001100111","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000100010","001000100010","001100100010","010101000100","010101000100","010000110011","001000100001","001000100001","001000100001","001000100001","001000100010","010100110011","011101000100","100001000101","100001010101","010000110011","001000100001","001000100001","001000100001"),
		("011101100110","001100100010","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010000110100","010101000100","010000110011","001000100001","001000100001","001000100001","001000100001","001000010001","010100110011","011101000100","100001000101","100001010110","011000110100","001000100001","001000100001","001000100010"),
		("100001100111","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010101000100","001100110011","001000100001","001000100001","001000100001","001000010001","001000010001","010000100010","011100110100","011101000101","100001010110","011000110100","001000100001","001000100001","001000100001"),
		("100001100111","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010101000100","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","010100110011","011101000101","100001010101","010000110011","001000100001","001000010001","001000100001"),
		("100001111000","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110100","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","000100010001","001100100001","011000110011","011000110100","001100100010","001000100001","001000100001","001000100001"),
		("100101111001","011101010110","001100100010","001000100001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","010000110011","010000110100","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100001","001100100001","001000100001","001000100010","001100110011","001000100010"),
		("100110001001","011101010110","001100100010","001100100010","010000110011","010100110011","010100110011","010000110010","001000100001","001000010001","001000010001","001100110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010"),
		("100110001001","011101010110","001000100001","010000110011","011101010101","100101100110","100001010101","011101000100","001100100001","001000100001","001000100001","001100100010","010000110011","001100100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010"),
		("100110001001","100001111000","010000110011","010000110011","100001010101","100001000101","011101000100","011000110011","001100100001","001000010001","001000010001","001000100010","001100110011","001100100010","001000010001","001000100001","001000010001","001000010001","001000100001","001000100010","001000010001","000100010001","000100010001","001000010001","001000100001","001000100001","001100110011"),
		("100110001001","100110001001","100001111000","010101000100","011000110100","011000110011","011000110011","011000110011","001100100001","000100010001","001000010001","001000010001","001100100010","001100100010","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","000100010000","001000010001","001100110011","010000110011","010101000101","100001111000"),
		("100110001001","100010001001","100110001001","100001111000","011101000101","011000110011","011100110011","011000110011","001000100001","001000010001","001000010001","001000010001","001100110010","001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","000100010001","001100100010","100001110111","100110001001","100110001001","100110001001"),
		("100110001001","100010001001","100010001001","100010001001","100001111000","011000110011","011000110011","010000100010","001000010001","001000010001","001000010001","001000100010","001100110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001100100010","011101100111","100110001001","100110001001","100110001001"),
		("100010001001","100001111000","100001111000","100010001001","011101100111","001100100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000100001","001100110010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","010101000101","100110001001","100110001001","100110001001"),
		("100001111000","100001111000","100001111000","100001111000","010101000101","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001100110010","001000100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100001","010000110100","100001111001","100110001001","100110001001"),
		("100001111000","100001111000","100001111000","100001111000","010000110011","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001100110011","001100100010","001000010001","001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","001000100001","001000010001","010000110011","100001111000","100010001001","100010001001"),
		("100001110111","100001100111","100001110111","011101100111","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","001100100010","001000100010","001000010001","001000010001","001000010001","001000010001","001100110011","001000100001","000100010001","001000010001","001000010001","001100100010","011101100111","100001111000","100001111000"),
		("011001100110","011001100110","011101100110","011001010101","001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001100100010","011001010110","011101100111","011101100111"))
	-- 10
	,

		(	("101010011100","101010101100","101010101100","101010101100","101010101100","100110011011","100101110111","100101100101","100101100101","100001010100","011100110011","010000100001","010000100001","010000100001","010000100010","001100100001","001100010001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","010000100010"),
		("101110101100","101110101101","101110101100","101110101101","101010101100","100101111000","100101010101","011101000011","011101000011","011100110011","010100100010","001100100001","001100010001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","010000100001","010000100010"),
		("101110101100","101110101100","101110101100","101110101100","101010001001","100101100101","011101000011","010100100010","010100100010","010100100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100001","010000100010","010000100010","010000100010","010000100010","010000100001","001100100001","010000100010","010000100001"),
		("101110101101","101110101101","101110101101","101110101100","100101100110","100001010100","100001000011","011000110011","010100100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","010000100001","010000100010","010000100010","010100100010","010000100010","010000100001","010000100001","001100100001","001100100001","010000100001","001100100001"),
		("101010101100","101010011100","101010011011","100110001010","100101010101","011101000011","011101000011","010100110010","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100100001","010000100001","010000100010","001100100001","010000100001","010000100001","010000100001","001100100001","001100010001","001100100001","001100100001","001100100001"),
		("100110001010","100110001011","100110011011","100101111001","100101100110","011101000011","010100100010","010000100001","010000100001","010000100001","010000100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001"),
		("100110001011","100110011011","100110011011","100110001010","100101111001","100001100110","010100100010","010000100001","001100100001","010000100001","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100101100111","011100110011","010100100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100001","010000100010","001100100001","001100100001"),
		("100110011011","100110011011","100110011011","100110001010","100110001011","100110001001","100001000101","011000110010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100010","010000100010","010000100010","010100100010","010000100010","010000100010","010000100010","010000100010"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","100110001010","100101111000","011101000100","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010100100010","010100110011","010100110011","011000110011","011000110011","010100110011","010100110011","010100100010"),
		("100110011011","100110011011","100110011011","100110011011","100110001010","100110001010","100110001001","100101100111","011000110011","010100100010","010000100001","010000100001","001100100001","010000100001","010000100001","010000100010","010000100010","010100100010","011000110011","011000110100","011101000100","011101000101","011101000101","011101000101","011101000100","011000110011","010100110011"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100110001010","100101111001","011101000101","011000110011","010100110011","010000100010","010000100010","010100100010","010100110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010101","100001010101","100001010110","100001010110","100001000101","011101000100","011000110011"),
		("100110001010","101010011011","101010011011","100110011011","100110001010","100001111001","100010001001","100101111001","100001010101","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110100","011000110100","011101000100","100001000101","100001010101","100001010110","100001010110","100001010110","100001010110","100001010110","011101000101","011000110011"),
		("101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001","100001111000","011101000101","011101000100","011101000100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","011101000101","011000110011"),
		("101010101100","101010101100","101010011100","101010011011","100010001001","100001111001","100001111001","100001100111","011101000100","011101000100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100101010111","011101000101","011000110100"),
		("101010101100","101110101100","101010101100","101010011011","100010001001","100001111001","100001111001","100001100111","011101000100","011101000100","011000110100","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110","100101010111","100001010101","011101000100"),
		("101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","100010001010","100001100111","011101000100","011001000100","011000110100","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001010110","100001010110","100001010111","100001010110","011101000100"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","100110001011","100110001010","100101100111","100001000101","011101000100","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010111","100001010110","011101000100"),
		("101010011011","101010011011","101010011011","101010011011","100110011011","100110011010","100110001001","100101100111","100001010101","011100110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010111","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100101100111","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110","100001010111","100001010111"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","100110011011","100110001001","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000101","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101010101100","101010011100","100110001001","100001100110","011000110011","010100100010","010100110010","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","101110101100","100110001010","100101111000","011101000101","011000100011","010100100010","010100100010","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000101","100001010110","100001010110","100001010111"),
		("101110111101","101110111101","101110111101","101110101101","101110111101","101010101100","100110001010","100010001001","100001010110","011000110011","010100100010","010100100010","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","011000110011","011101000100","100001000101","100001010110","100001010111"),
		("101110111101","101110111101","101110111101","101110101101","101110101101","101010011100","100110001010","100010001001","100101100111","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000100","100001000101","100001010110","100101010111"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010101100","100110001010","100110001001","100101100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","011000110011","011000110100","011101000100","011101000100","100001000101","100001010110","100101010111"),
		("101110101101","101110101101","101110101101","101110101101","101110111101","101010011011","100110001010","100110001001","100001010110","011000110100","011100110100","011100110100","011101000100","011101000100","011101000100","011000110011","011000110011","011000110011","011000110010","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110","100001010111"),
		("101110111101","101110101101","101110101101","101110101101","101110101101","101010011011","100110001010","100110001001","100001010101","011000110100","011101000100","011101000100","100001010110","100001010110","100001000101","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010011100","100110001010","100110001001","100001010110","011101000100","100001010101","011101000101","100001010110","100001010111","100001010110","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101110111101","101010011011","100110001010","100110001010","100001100111","100001010101","011101000101","011101000101","100001010110","100001010111","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100110001010","100101111000","011101000101","011000110100","011101000101","100001000101","100001000101","100001010110","011101000100","011000110010","010100100010","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","100110001001","011101000100","011000110011","011100110100","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010011010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001010101","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","101010011011","101010011011","011101010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010101","100001010110","100001010110","100001010110"),
		("101110111101","101110111110","101110111110","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","100001111000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010101","100001010101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011100","101110101101","101010011010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001010101","100001010110","100001010110"),
		("101110111101","101110101101","101110101101","101110101100","101010011011","100110011011","100110011011","101010011011","101010101100","101010101100","100001101000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110010","011000110011","011000110011","011100110100","100001000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111101","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","101010101100","101110101100","101110101100","101010011011","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001010101","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","100110011011","100110011011","100110011011","101010101100","101010101100","101010101100","101010101100","100101111000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","100001000101","100001010101"),
		("101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","100110011011","101010101100","101110101100","101010101100","101010011100","100110001010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","011101000100","011101000100","011101000101","100001000101","100001000101"),
		("101110111101","101110111101","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","101110101101","100001111001","010100110100","010101000100","010101000100","010101000100","010101000100","011001000100","011101100110","011101000101","011000110011","011000110100","011101000100","100001000101","100001000101","100001000101","100001000101","100001000101","100001000101"),
		("101110111101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011011","101110101101","101110101101","011101100111","010000110011","010000110011","010001000100","010101000100","010101000101","010101000101","011101100111","011101010110","011000110100","011101000100","011101000100","011101000101","011101000101","011101000100","011101000100","011101000100","011101010101"),
		("101110101101","101110111101","101110111101","101010011011","100110011011","100110011011","101010011100","101110101101","101110101100","100001111000","011001000101","010001000100","010000110011","010000110011","001100110011","010101000100","010101010101","010101000100","011101000100","011101000100","011101000100","011101000100","011000110100","011000110011","011000110011","011101000100","100001010101"),
		("101110111101","101110111101","101110111101","101010011011","100110011011","100110011011","101010101100","101110101101","101110101100","100001111001","010101000100","010101000100","010101000100","010000110011","010000110011","010101000100","010101010101","010101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","100001010101"),
		("101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010101100","101110101101","101110101101","100001111001","010100110100","010001000100","010101000100","010101000100","010000110100","010101000100","011001010101","011001010101","011101000100","011000110011","011000110010","011000110010","011000110011","011000110011","011000110011","011000110011","011101000101"),
		("101010101100","101110101101","101010011100","100110011011","100110011011","100110011011","101010101100","101010101100","101010101100","100001111000","010000110011","010000110011","010000110011","010000110011","010000110100","010101000101","011001010101","011001010101","011000110011","011000110010","010100100010","011000100010","011000110011","011000110011","011000110011","011000110011","011100110100"),
		("101010011100","101010101100","100110011011","100010001010","100110001010","100110001010","100110011011","101010011011","100110011011","011101100111","010000110011","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010101","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100110010"),
		("100110001010","100110001010","100001111001","100001111000","100001111001","100001111001","100010001010","100110001010","100110001010","011001010110","001100110011","001100100011","001100100011","001100110011","001100110011","010000110100","010101000100","010101000100","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010"))
	-- 11
	,

		(	("101010011100","101010101100","101010101100","101010101100","101010101100","101010011011","101010011011","100110011010","100110011011","100010001001","100001100111","100001010101","011000110011","010100100010","010100110010","011000110011","011000110011","011000110010","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011000110011","010100110010"),
		("101110101100","101110101101","101110101100","101110101101","101010101100","101010101100","101010101100","101010011011","101010011011","100110001001","100101100111","100001000101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000101","011101000101","011101000101","011101000101","011101000100","011000110011"),
		("101110101100","101110101100","101110101100","101110101100","101010101100","101010101100","101010011100","101010011011","101010011011","100101111001","100001010110","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001000101","100001000101","011101000101","011000110011"),
		("101110101101","101110101101","101110101101","101110101101","101110101101","101110101100","101010101100","101010101100","101010011011","100101111000","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001010110","011101000101","011000110011"),
		("101010101100","101010011100","101010011011","101010011100","101010011011","101010011011","100110001010","100110001010","100110001010","100101111000","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000100","100001000101","100001010110","100001000101","011000110100"),
		("100110001010","100110001011","100110011011","100110001011","100110001010","100110001010","100010001010","100001111001","100001111001","100001111001","100001010110","011100110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001000101","011100110100"),
		("100110001011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001","100101111000","100001010101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","011101000100"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100101111000","100001000101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001010110","100001010110","100001000101"),
		("100110011011","100110011011","100110011011","100110001010","101010011011","101010011011","100110011011","100110011011","100110001001","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","101010011011","101010011011","100110001010","100001111001","011101010101","011000100010","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001010","100110001010","101010011011","101010011011","100010001001","100001101000","011000110011","010100100010","011000110011","011000110011","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110010","011000110011","011101000100","011101000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100110001010","101010011011","100010001010","100001111001","011101010101","010100100010","010100110011","011000110011","011000110011","011000110011","010100110011","010000100010","010100100010","010100100010","010100110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110"),
		("100110001010","101010011011","101010011100","100110011011","100110001010","100001111001","100010001001","100110001010","100010001010","100010001001","100001100111","011000110100","011000110100","011000110011","011000110011","011000110100","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000101","100001010110","100001010110"),
		("101010011011","101010011011","101010011011","101010011100","100010001001","100001111001","100001111001","100010001001","100010001010","100010001001","100101100111","100001010101","011101000100","011000110011","011000110100","011000110100","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100001010110","100001010110"),
		("101010101100","101010101100","101010011100","101010011011","100010001001","100001111001","100001111001","100010001001","100010001010","100101111001","100101100111","100001010101","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101010101100","101110101100","101010101100","101010011011","100010001001","100001111001","100001111001","100010001001","100010001010","100101111000","100001010110","011000110100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","100010001001","100010001001","100010001010","100101110111","011101000100","011101000101","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001010101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011011","101010011011","100110001011","100110001010","100010001001","100010001001","100001010101","011100110100","100001000101","100001010110","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101010011100","101010011100","101010011011","101010011011","100110011011","100110011010","100110001001","100001111001","100001111001","011101010101","011000110100","011100110100","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","100001000101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111001","100001100111","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001000110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111001","100001111000","100001010101","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","011101000100","100001000101","100001000101","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101010101100","101010011100","100110001010","100001111001","100001111001","100001111001","100101100111","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","101110101100","100110001010","100001111001","100010001010","100110001010","100101100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110111101","101010101100","100110001010","100001111001","100010001001","100110011010","100101100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110101101","101010011100","100110001010","100010001001","100010001010","101010011011","100110001001","011101000100","011000110011","011000110011","011000110010","011000110010","011000110010","010100100010","010100100010","011000110011","011000110011","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010101100","100110001010","100110001010","100110001010","101010011011","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","011000110010","011000110011","011000110011","011000110100","011101000100","011101000100","100001000101","100001000101","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001001","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","100001000101","100001000101","100001000101","100001000101"),
		("101110111101","101110101101","101110101101","101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010001010","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011100110100","011101000100","011101000100","100001000101","100001000101"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010011100","100110001010","100110001010","100110011011","101010101100","101010101100","101010011011","100001100110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011000110100","011101000100","011101000100","011101000100","011101000101","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101110111101","101010011011","100110001010","100110001010","101010011011","101010101100","101010101100","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000101","011101000101","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100110001010","101010011011","101010011100","101010011100","101010101100","100101111000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101010101100","101010011011","100001100111","011000110100","011000110011","011000100010","011000110011","011000110011","011000110011","011000110100","011101000100","011100110100","011000110011","011000110011","011100110100","011101000100"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010101100","101110101101","101110101100","101010101100","101010101100","101110101100","101010011011","100101111000","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","101010011011","101010101100","101110101100","101010101100","101010101100","101010101100","101010101100","101110101100","101010101100","100001111000","011101000100","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110"),
		("101110111101","101110111110","101110111110","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","101110101101","101110101101","101110101100","101110101100","101110101101","101010101100","100001101000","011000110011","100001010101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011011","101110101101","101110101101","101110101101","101110101100","101010101100","101010011011","011101100110","011000110011","011000110011","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101"),
		("101110111101","101110101101","101110101101","101110101100","101010011011","100110011011","100110011011","101010011011","101110101100","101010011100","101010011010","100001111000","011101010110","011001000100","011000110011","011000110011","011101000100","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100"),
		("101110111101","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","101010011011","100110001010","011101100110","011001000100","011000110011","011000110011","011000110011","011000110011","011000110011","100001010110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100001111000","011001010110","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","100101100110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101110111101","101110101101","100110011011","100001111000","011001010101","010100110011","010100110011","010100110011","010100110011","010000100010","010000100010","010000100010","010100100010","010100100011","011001000100","100101100111","011101010110","010100110011","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101010011100","100001111000","011001010101","010100110011","010100100010","010000100010","010000100010","010101000100","010100110011","010000110011","010000110011","010101000100","010101000100","010101000100","011101100110","100101111000","011101100110","010100110011","010000100001","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("100110001001","011001010101","011000110011","010100110011","010000100010","010000100001","001100100001","001100100001","010000110011","010000110011","010000110011","010000110011","010000110100","010101000100","010101000101","011101100110","011101100111","011101100110","011001000100","010000100001","010000100010","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("011001000100","010100110011","010100100010","010000100010","001100100001","001000100001","001000010001","001000010001","010000100010","010101000101","010101000100","010000110011","010000110011","001100110011","010000110100","011001010110","010101000100","011101100110","011001010101","010000100010","010000100001","010100100010","010100110011","011000110011","011000110011","011000110011","011000110011"),
		("010100110011","010000100010","001100100001","001000100001","001000010001","001000010001","001000010001","001000010001","001100110010","010101000100","010000110100","010001000100","010000110100","010000110011","010000110011","011001010101","010101000101","011101100110","011101100110","010100110011","010000100001","010000100001","010100100010","011000110011","011000110011","011000110011","011000110011"),
		("010000100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100100010","010100110100","010000110011","010000110100","010000110100","010000110100","010001000100","011001010110","011001010101","011101100111","100001111001","011101100111","010100100010","010100100010","010100100010","011000110011","011000110011","011000110011","011000110011"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100110010","010100110100","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010110","011101100111","100001111000","100001111001","011001000100","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","010000110011","001100110011","001100110011","001100110011","010000110011","010000110100","011001010101","011001010101","011001010110","011101100110","100001111000","011101100111","010100110010","010100100010","010100100010","010100100010","010100100010","010100110010"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","001100110011","001100100010","001100100010","001100100010","001100100011","010000110011","010101000100","010101000100","011001010101","010101010101","011101100110","011101100111","010100110100","010100100010","010100100010","010100100010","010100100010","010100100010"))
	-- 12
	,

		(	("101010011100","101010101100","101010101100","101010101100","101010101100","101010011011","101010011011","100110011010","100110011011","100010001001","100001100111","100001010101","011000110011","010100100010","010100110010","011000110011","011000110011","011000110010","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011000110011","010100110010"),
		("101110101100","101110101101","101110101100","101110101101","101010101100","101010101100","101010101100","101010011011","101010011011","100110001001","100101100111","100001000101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000101","011101000101","011101000101","011101000101","011101000100","011000110011"),
		("101110101100","101110101100","101110101100","101110101100","101010101100","101010101100","101010011100","101010011011","101010011011","100101111001","100001010110","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001000101","100001000101","011101000101","011000110011"),
		("101110101101","101110101101","101110101101","101110101101","101110101101","101110101100","101010101100","101010101100","101010011011","100101111000","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001010110","011101000101","011000110011"),
		("101010101100","101010011100","101010011011","101010011100","101010011011","101010011011","100110001010","100110001010","100110001010","100101111000","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000100","100001000101","100001010110","100001000101","011000110100"),
		("100110001010","100110001011","100110011011","100110001011","100110001010","100110001010","100010001010","100001111001","100001111001","100001111001","100001010110","011100110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001000101","011100110100"),
		("100110001011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100001111001","100001111001","100101111000","100001010101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","011101000100"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100101111000","100001000101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001010110","100001010110","100001000101"),
		("100110011011","100110011011","100110011011","100110001010","101010011011","101010011011","100110011011","100110011011","100110001001","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","101010011011","101010011011","100110001010","100001111001","011101010101","011000100010","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001010","100110001010","101010011011","101010011011","100010001001","100001101000","011000110011","010100100010","011000110011","011000110011","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110010","011000110011","011101000100","011101000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100110001010","101010011011","100010001010","100001111001","011101010101","010100100010","010100110011","011000110011","011000110011","011000110011","010100110011","010000100010","010100100010","010100100010","010100110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110"),
		("100110001010","101010011011","101010011100","100110011011","100110001010","100001111001","100010001001","100110001010","100010001010","100010001001","100001100111","011000110100","011000110100","011000110011","011000110011","011000110100","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000101","100001010110","100001010110"),
		("101010011011","101010011011","101010011011","101010011100","100010001001","100001111001","100001111001","100010001001","100010001010","100010001001","100101100111","100001010101","011101000100","011000110011","011000110100","011000110100","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100001010110","100001010110"),
		("101010101100","101010101100","101010011100","101010011011","100010001001","100001111001","100001111001","100010001001","100010001010","100101111001","100101100111","100001010101","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101010101100","101110101100","101010101100","101010011011","100010001001","100001111001","100001111001","100010001001","100010001010","100101111000","100001010110","011000110100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","100010001001","100010001001","100010001010","100101110111","011101000100","011101000101","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001010101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011011","101010011011","100110001011","100110001010","100010001001","100010001001","100001010101","011100110100","100001000101","100001010110","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101010011100","101010011100","101010011011","101010011011","100110011011","100110011010","100110001001","100001111001","100001111001","011101010101","011000110100","011100110100","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","100001000101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111001","100001100111","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001000110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111001","100001111000","100001010101","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","011101000100","100001000101","100001000101","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101010101100","101010011100","100110001010","100001111001","100001111001","100001111001","100101100111","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","101110101100","100110001010","100001111001","100010001010","100110001010","100101100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110111101","101010101100","100110001010","100001111001","100010001001","100110011010","100101100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110101101","101010011100","100110001010","100010001001","100010001010","101010011011","100110001001","011101000100","011000110011","011000110011","011000110010","011000110010","011000110010","010100100010","010100100010","011000110011","011000110011","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010101100","100110001010","100110001010","100110001010","101010011011","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","011000110010","011000110011","011000110011","011000110100","011101000100","011101000100","100001000101","100001000101","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101110111101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","100110001001","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","100001000101","100001000101","100001000101","100001000101"),
		("101110111101","101110101101","101110101101","101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010001010","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011100110100","011101000100","011101000100","100001000101","100001000101"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010011100","100110001010","100110001010","100110011011","101010101100","101010101100","101010011011","100001100110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011000110100","011101000100","011101000100","011101000100","011101000101","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101110111101","101010011011","100110001010","100110001010","101010011011","101010101100","101010101100","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000101","011101000101","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100110001010","101010011011","101010011100","101010011100","101010101100","100101111000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010011100","101110101101","101110101100","101010101100","101010011011","100001100111","011000110100","011000110011","011000100010","011000110011","011000110011","011000110011","011000110100","011101000100","011100110100","011000110011","011000110011","011100110100","011101000100"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010101100","101110101101","101110101100","101010101100","101010101100","101110101100","101010011011","100101111000","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","101010011011","101010101100","101110101100","101010101100","101010101100","101010101100","101010101100","101110101100","101010101100","100001111000","011101000100","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110"),
		("101110111101","101110111110","101110111110","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","101110101101","101110101101","101110101100","101110101100","101110101101","101010101100","100001101000","011000110011","100001010101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011011","101110101101","101110101101","101110101101","101110101100","101010101100","101010011011","011101100110","011000110011","011000110011","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101"),
		("101110111101","101110101101","101110101101","101110101100","101010011011","100110011011","100110011011","101010011011","101110101100","101010011100","101010011010","100001111000","011101010110","011001000100","011000110011","011000110011","011101000100","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100"),
		("101110111101","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","101010011011","100110001010","011101100110","011001000100","011000110011","011000110011","011000110011","011000110011","011000110011","100001010110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100001111000","011001010110","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","100101100110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101110111101","101110101101","100110011011","100001111000","011001010101","010100110011","010100110011","010100110011","010100110011","010000100010","010000100010","010000100010","010100100010","010100100011","011001000100","100101100111","011101010110","010100110011","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111101","101010011100","100001111000","011001010101","010100110011","010100100010","010000100010","010000100010","010101000100","010100110011","010000110011","010000110011","010101000100","010101000100","010101000100","011101100110","100101111000","011101100110","010100110011","010000100001","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("100110001001","011001010101","011000110011","010100110011","010000100010","010000100001","001100100001","001100100001","010000110011","010000110011","010000110011","010000110011","010000110100","010101000100","010101000101","011101100110","011101100111","011101100110","011001000100","010000100001","010000100010","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("011001000100","010100110011","010100100010","010000100010","001100100001","001000100001","001000010001","001000010001","010000100010","010101000101","010101000100","010000110011","010000110011","001100110011","010000110100","011001010110","010101000100","011101100110","011001010101","010000100010","010000100001","010100100010","010100110011","011000110011","011000110011","011000110011","011000110011"),
		("010100110011","010000100010","001100100001","001000100001","001000010001","001000010001","001000010001","001000010001","001100110010","010101000100","010000110100","010001000100","010000110100","010000110011","010000110011","011001010101","010101000101","011101100110","011101100110","010100110011","010000100001","010000100001","010100100010","011000110011","011000110011","011000110011","011000110011"),
		("010000100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100100010","010100110100","010000110011","010000110100","010000110100","010000110100","010001000100","011001010110","011001010101","011101100111","100001111001","011101100111","010100100010","010100100010","010100100010","011000110011","011000110011","011000110011","011000110011"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100110010","010100110100","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010110","011101100111","100001111000","100001111001","011001000100","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","010000110011","001100110011","001100110011","001100110011","010000110011","010000110100","011001010101","011001010101","011001010110","011101100110","100001111000","011101100111","010100110010","010100100010","010100100010","010100100010","010100100010","010100110010"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001100100010","001100110011","001100100010","001100100010","001100100010","001100100011","010000110011","010101000100","010101000100","011001010101","010101010101","011101100110","011101100111","010100110100","010100100010","010100100010","010100100010","010100100010","010100100010"))
	-- 13
	,

		(	("101010011100","101010101100","101010101100","101010101100","101010101100","101010011011","101010011011","100110011010","100110011011","100001111001","100001100111","011101000100","011000110011","010100110010","010100110011","011000110011","011000110011","011000110010","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011100110100","010100100010","010100100010"),
		("101110101100","101110101101","101110101100","101110101101","101010101100","101010101100","101010101100","101010011011","101010011011","100110001001","100101100111","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000101","011101000101","011101000101","011101000100","011000110011","011000110010"),
		("101110101100","101110101100","101110101100","101110101100","101010101100","101010101100","101010011100","101010011011","101010011011","100101111001","100001010110","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","100001000101","100001000101","100001000101","011000110011","010100100010"),
		("101110101101","101110101101","101110101101","101110101101","101110101101","101110101100","101010101100","101010101100","101010011011","100101111000","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001000101","100001000101","011101000101","011000110011","010100100010"),
		("101010101100","101010011100","101010011011","101010011100","101010011011","101010011011","100110001010","100110001010","100110001010","100101110111","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","100001000101","100001000101","100001000101","011000110011","011000110011"),
		("100110001010","100110001011","100110011011","100110001011","100110001010","100110001010","100010001010","100001111001","100001111001","100101100111","100001000101","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001010110","011000110011","011000110011"),
		("100110001011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001100110","011101000100","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100001000101","100001000101","100001010110","011100110100","011000110011"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100001111001","100001010110","011100110100","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","100001000101","100001000101","100001000101","100001010110","011101000101","011000110011"),
		("100110011011","100110011011","100110011011","100110001010","101010011011","101010011011","100110011011","100110011011","100101111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","100001000101","100001000101","100001000101","100001000101","100001010110","100001010110","011101000100"),
		("100110011011","100110011011","100110011011","100110011011","100110011011","101010011011","101010011011","100110001010","011101010101","010100100010","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","011101000100","100001000101","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001010","100110001010","101010011011","101010011011","100001100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100110010","011000110011","010100110010","010100100010","011000110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100110001010","101010011011","100101111000","011000110011","010100100010","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010100100010","010100100010","010100100010","011000110011","011000110100","011101000101","100001010110","100001010110","100001010110","100001010110"),
		("100110001010","101010011011","101010011100","100110011011","100110001010","100001111001","100010001001","100110001010","100110001001","011101000101","011001000100","011101000100","011000110011","011000110011","011000110100","011000110011","010000100010","010100100010","010000100010","010100100010","010100110010","011000110011","011101000100","100001010110","100001010110","100001010110","100001010110"),
		("101010011011","101010011011","101010011011","101010011100","100010001001","100001111001","100001111001","100010001001","100010001010","100101111000","100001010101","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110"),
		("101010101100","101010101100","101010011100","101010011011","100010001001","100001111001","100001111001","100010001001","100110001010","100001010110","011100110011","011000110011","011000110100","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110100","011100110100","011101000101","100001010110","100001010110","100001010110","100001010110"),
		("101010101100","101110101100","101010101100","101010011011","100010001001","100001111001","100001111001","100010001010","100001101000","011101000100","011101000100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","100010001010","100001111000","011101000101","011101000101","100001010110","100001000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001000101","100001010101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011011","101010011011","100110001011","100110001010","100001100111","011100110100","011101000101","100001000101","100001000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","100001000101","100001010110","100001010110"),
		("101010011100","101010011100","101010011011","101010011011","100110011011","100110011010","100110001010","100001111000","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","100001000101","100001000101","100001000101","100001010110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","100110001001","100001111001","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","100001000101","100001000101","100001000110","100001010110"),
		("101010101100","101010101100","101010101100","101010011100","101010011011","100110011011","100110001001","100001111001","100001100111","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001000101","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101010101100","101010011100","100110001010","100001111001","100101100111","100001010110","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","101110101100","100110001010","100010001001","100101111000","100001010101","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110111101","101010101100","100110001010","100010001001","100001111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001000110","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101110101101","101110101101","101010011100","100110001010","100010001001","100001111001","011000110100","011000110011","010100100010","011000110011","011000110011","011000110010","011000110010","011000110010","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001000101","100001010110","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010101100","100110001010","100110001010","100010001001","100001010110","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110010","011000110011","011101000100","011101000100","011101000100","011101000100","011101000101","100001000101","100001000101","100001010110"),
		("101110101101","101110101101","101110101101","101110101101","101110111101","101010011011","100110001010","100110001010","100110001010","100110001001","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","100001000101","100001000101","100001000101","100001000101"),
		("101110111101","101110101101","101110101101","101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","101010011011","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001000101"),
		("101110111110","101110111110","101110111110","101110111110","101110111110","101010011100","100110001010","100110001010","100110011011","101010101100","100101100111","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011000110100","011101000100","011000110100","011101000100","011101000100","011101000100","011101000101","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101110111101","101010011011","100110001010","100110001010","101010011011","101010101100","100101111000","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000100","011101000101"),
		("101110111101","101110111101","101110111101","101110111101","101110101101","100110011011","100110001010","100110001010","101010011011","101010011100","100101100111","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000101","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010011100","101110101101","101010011010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001000110"),
		("101110111101","101110111101","101110111101","101110111110","101110101101","100110011011","100110011011","100110011011","101010101100","101110101101","101110101100","100110001010","011101010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011100110100","011101000100","011101000101","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110011011","100110011011","101010011011","101010101100","101110101100","101010101100","101010101100","101010011100","101010011010","100001100111","011101000100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001010110"),
		("101110111101","101110111101","101110111110","101110111110","101010101100","100110011011","100110011011","101010011011","101110101100","101110101101","101110101101","101110101100","101110101101","101010011011","011101010101","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","100001000101","100001010110","100001010110","100001010110"),
		("101110111101","101110101101","101110111101","101110111101","101010011100","100110011011","100110011011","101010011011","101110101101","101110101101","101110101101","101010101100","100101111001","011001000100","011101000100","100001010110","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","100001000101","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101010101100","100110011011","100110011011","100110011011","101010011100","101010101100","101010011011","100110001010","011101010110","011000110011","011000110011","100001010101","100001000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","100001000101","100001010110","100001010110","100001010110"),
		("101110101101","101110101100","101110101101","101110101100","100110001011","100110001010","100110001001","100001111000","011101100110","011001000100","011000110011","011000110011","011000110011","011001000100","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010101","100001010110"),
		("101110111101","101110101101","101110101101","101010011010","011101100111","011001000101","011000110100","010100110011","010100110011","010100100011","010100110011","010100110011","010100110011","100001010101","100001010101","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101"),
		("101010011011","100001111000","011101010110","011000110100","010100110011","010000100010","010000100010","010000100010","010000100010","010100110010","010000100010","010100110011","010100110011","100101100110","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100"),
		("011001000100","011000110011","010100100010","010000100010","010000100010","001100100001","001100100001","001100100001","001100100001","011001000100","010000100010","010000110011","010100110100","011001000101","011001000101","011001000100","011101010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100"),
		("010100110011","010000100010","010000100001","001100100001","001000100001","001000010001","001100100001","001100100001","001100100001","010000110011","010000110011","010000110011","010001000100","010101000100","010101000100","010101010101","011101100111","011001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100"),
		("010000100010","001100100001","001000010001","001000010001","001000010001","001000100001","001000010001","001000010001","001000010001","010000110011","010101000100","010000110011","010000110011","001100110011","001100110011","010101000101","010101000101","010100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010100110100","010000110100","010000110100","010000110100","010000110011","010000110011","010101000100","010101000101","010100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","010000110011","010000110011","010000110100","010000110011","010101000100","011001010101","010101000100","011000110011","011000110011","011000110010","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","010000110011","010000110011","010000110011","010000110011","010101000101","011001010101","010101000100","010100100010","011000110011","011000110011","011000100010","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010000110011","010000110011","001100110011","001100110011","001100110011","010000110011","010101000100","011001010101","010101000100","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100110010"),
		("000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000010001","010000110011","001100100010","001100100010","001100100010","001100100011","001100110011","010000110100","010101000100","010000110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010"))
	-- 14
	,

		(	("101010011100","101010101100","100101111000","011101000100","010100100010","010000100001","010000100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100010001","001100010001"),
		("101110101100","101010101100","100001100111","011000110010","010100100010","010000100001","010000100001","001100100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("101110101100","101010011011","100001100111","011001000100","010100100010","010100100010","010000100001","010000100001","001100100001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("101110101101","101110101101","101010011011","100101111000","011000110011","010100100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("101010101100","101010011100","101010011011","100001111000","011101000100","010100110010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100010","001100100001","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001"),
		("100110001010","100110001010","100110001010","100001111000","011101000101","010100100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100010","010100100010","010100100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001"),
		("100110001011","100110011011","100110001010","100001111001","100001010110","011000110010","010000100001","001100100001","001100100001","010000100001","010000100010","010000100010","010100100010","011000110011","011000110011","011000110011","011100110011","011100110100","011000110011","010100110011","010100100010","010000100010","010000100001","010000100001","001100100001","001100100001","001100100001"),
		("100110011011","100110011011","100110011011","100110001010","100101111001","011101000101","010100100010","010000100010","010100100010","011000110011","011000110011","011000110011","011000110100","011000110011","011100110100","011101000100","011101000100","011101000100","011101000100","011000110011","011000110011","010100100010","010100100010","010000100010","010000100010","010000100010","010000100001"),
		("100110011011","100110011011","100110011011","100110001010","100110001010","100101100111","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","011101000101","011101000101","011101000101","011101000100","011100110100","011000110011","010100100010","010100100010","010000100010","010000100010","010000100001"),
		("100110011011","100110011011","100110001011","100110001010","100110001010","100101100110","011101000100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000101","100001000101","100001000101","100001000101","100001000101","011101000101","011000110011","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001"),
		("100110011011","100110011011","100110001010","100110001010","100101111000","100001010101","011101000100","011101000100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100001000101","100001000101","100001000101","100001010110","011101000101","011000110011","011000110011","010100100010","010000100010","010000100010","010000100010","010000100001"),
		("100110011011","100110011011","100110011011","100110001010","100101110111","100001010101","011101000100","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000101","100001010110","100001010110","100001000101","011000110011","011000110011","010100100010","010000100010","010000100010","010000100010","001100100001"),
		("100110001010","101010011011","101010011100","100110011011","100101110111","100001010101","011101000100","011100110011","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001010110","100001010110","100001000101","011100110100","011000110011","010100100010","010000100010","010000100010","010000100010","001100100001"),
		("101010011011","101010011011","101010011011","101010011011","100101111000","100001010101","011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110100","011000110011","011000110100","011000110100","100001000101","100001010110","100001010110","100001010110","011101000100","011000110011","010100110010","010000100010","010000100001","010000100010","010000100010"),
		("101010101100","101010101100","101010011100","101010011011","100101111000","011101000100","011100110011","011100110011","011000110011","011000110011","011000110011","011000110011","011000110100","011000110100","011000110100","011100110100","100001000101","100001010110","100001010110","100001010110","100001000101","011100110100","010100100010","010000100010","010100100010","010000100010","010000100010"),
		("101010101100","101110101100","101010101100","101010011011","100101100111","011101000100","011000110011","011100110011","011000110011","011000110100","011000110100","011000110011","011000110100","011000110100","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","011101000101","011000110011","010100100010","010100100010","010100100010","010100100010"),
		("101010011100","101010011100","101010101100","101010011011","100001100110","011100110011","011000110011","011000110011","011000110011","011000110011","010100110010","010100100010","010100110010","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001000101","011000110011","010100110011","010100110011","010100110011"),
		("101010101100","101010101100","101010101100","100110001010","011101000100","011000110011","011000110011","011000110011","011000110010","010100100010","010100100010","010100100010","010100100010","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","011101000101","011000110011","011000110011","011000110011"),
		("101010011100","101010011100","101010011100","100110001010","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100110010","011000110011","011000110011","011000110011","011101000101","100001000101","100001010110","100001010110","100001010110","100001010111","100001000101","011000110100","011000110011","011000110011"),
		("101010101100","101010101100","101010101100","101010011100","100001100111","011000110011","010100110010","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010100100010","011000110010","011000110011","011000110011","011000110100","100001000101","100001010110","100001010110","100001010110","100001010111","100001010110","011101000100","011000110011","011000110011"),
		("101010101100","101010101100","101010101100","101010011100","100110001001","011000110100","011000110100","011000110011","011000110011","011000110100","011000110011","010100100010","010000100010","010100100010","010100110011","011000110011","011000110011","011000110011","011101000100","100001010110","100001010110","100001010110","100001010111","100001010110","011101000100","011000110100","011000110100"),
		("101110101101","101110101101","101110101101","101110101101","101010011011","100101100111","100001000101","011000110011","011000110011","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","100001000101","100001010110","100001010110","100001010110","100001010111","100001010111","100001000101","011101000100","011101000100"),
		("101110111110","101110111110","101110111110","101110111101","101110101101","100101111000","011100110011","011000110011","011000110011","011100110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","100101010111","100001010110","100001000101"),
		("101110111101","101110111101","101110111101","101110111101","101010011100","100001010101","011101000100","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","100101010111","100101010111","100101100111"),
		("101110111101","101110111101","101110111101","101110101101","100001100111","011101000100","100001010110","011101000101","011000110100","011000110011","011000110011","011000110010","011000110011","011000110011","011000110010","011000110011","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100101010111","100101010111","100101010111"),
		("101110111110","101110111110","101110111110","101010011011","011101000100","011101000101","100001000101","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100101010111","100101010111","100101010111"),
		("101110101101","101110101101","101110101101","101010011011","100001010110","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000101","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100101010111","100101010111","100001010110"),
		("101110111101","101110101101","101110101101","101110101101","100110001001","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001000101","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","100101010111","100001010110"),
		("101110111110","101110111110","101110111110","101110111110","101010001010","011101000101","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000101","011101000101","100001000101","100001010110","100001010110","100001010110","100101010111","100101010111","100001010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101010011011","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110","100101010111","100101010111","100001010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100101100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010111","100101010111","100101010111","100001010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101100","100001100111","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010111","100101010111","100101010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111110","101110101100","100001100111","011000110011","011000110011","011000110010","011000110010","011000100010","010100100010","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010111","100001010111","100001010110"),
		("101110111101","101110111101","101110111101","101110111101","101010101100","100110001001","011101000100","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000101","100001000101","100001000110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111110","101110111110","101010101100","100110001010","100001100111","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110101101","101110111101","101110111101","101010011100","100110011011","100101111001","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","100001000101","100001000101","100001000101","100001010110","100001000101","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","101010101100","100110011011","100110011011","100110001010","100001100110","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001000101","100001000101","100001000101","100001000101","100001010110","100001010110","100001010110"),
		("101110101101","101110101100","101110101101","101110101100","100110001010","100110001010","100110001010","100101111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110011","011101000100","011101000100","011101000100","011101000100","100001000101","011101000101","100001000101","100001000101","100001010110","100001010110","100001010110","100001010101"),
		("101110101101","101110101101","101110101101","101110101100","100110001010","100110001010","100110001010","100101111001","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001000101"),
		("101110101101","101110101100","101110101101","101010101100","100110001010","100110001010","100110001010","101010011011","011101010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010101","100001010110","100001010110","100001000101"),
		("101110111101","101110111101","101110111110","101010011100","100110001011","100110001010","100110011011","101010101100","100101111000","010100100010","010100110011","010100110100","010100110100","010101000100","010101000100","011101010110","011101000101","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110111101","101110111101","101010011011","100110001011","100110001010","101010011011","101110101100","100001101000","010000100010","010000110011","010000110100","010001000100","010101000100","010101000101","011101100111","011001010101","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","101110101101","100110011011","100110011011","100110001010","101010011011","101010101100","100101111001","011001000101","010000110100","010000110011","001100110011","001100110011","010101000100","011001010101","010100110100","011000110011","011000110011","011000110011","011101000100","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110111110","101110101101","100110011011","100110011011","100110001010","101010011011","101110101100","100001111001","010100110100","010000110100","010000110100","010000110011","010000110011","010000110100","011001010101","010101000100","011000110011","011000110011","011000110011","011101000100","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110111101","101010101100","100110001010","100110001010","100110001010","101010011011","101010011010","011101100111","010000110011","010000110100","010000110100","010101000100","010000110011","010101000100","011001010110","010101000101","011000110011","011000110011","011000110011","011100110100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","100110001010","100001111001","100001111001","011101100111","011101010110","011001000100","010101000100","010000110011","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010101","011000110011","011000110011","011000110010","011000110011","011101000100","011101000100","011101000101","100001000101","100001000101","100001010110"),
		("100110001010","100110001001","011101100110","011001000100","010100110011","010000100010","010000100001","001100100001","010000110011","010000110011","001100110011","001100110011","001100110011","010000110011","010101000100","011001010101","011001000101","010100110011","010100100010","010100100010","010100110010","011000110011","011000110011","011000110100","011101000100","011101000100","100001000101"),
		("011001000101","010100110011","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000110011","001100100011","001100100010","001100100010","001100100010","001100110011","010000110011","010101000100","010101000100","010100100010","010100100010","010100100010","010100100010","010100100010","010100110010","011000110011","011000110011","011000110100","011101000100"))
	-- 15
	,

		(	("101010011100","101010101100","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111000","100001111001","100110001010","100110001010","100110001001","100001111001","100001111000","100010001001","100010001001","100110001010","100110001010","100110001010","100110011010","100110001010","100001111001","100001111001"),
		("101110101100","101110101100","101010101100","101110101100","101010101100","101010101100","101010101100","101010011100","101010101100","100110001010","100001111001","100001111001","100110001010","101010011011","100110001011","100110001010","100110001010","100110001010","101010011010","100110011011","101010011011","101010011011","101010011011","101010011011","100110001010","100010001001","100010001010"),
		("101110101100","101010101100","101010101100","101010101100","101010101100","101010011100","101010011100","101010011011","101010011011","100110001001","100001111001","100001111000","100001100111","100001100111","100001111000","100101111000","100101111001","100110001001","100110001010","100110011010","101010011011","101010011011","101010011011","101010011011","100110001010","100010001010","100010001010"),
		("101110101101","101110101101","101110101100","101110101101","101010101100","101010101100","101010011010","100110001001","100101100111","100001010101","011101000100","011000110011","011000110011","011000110010","011000110011","011000110011","011101000100","011101000100","100001010110","100101111000","100110001001","100110001001","100101111001","100110001001","100110001010","100010001001","100010001010"),
		("101010011100","101010011011","101010011011","101010011011","100110001001","100101100110","100001010100","011101000011","100001000011","011101000011","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","011000110011","011100110011","011101000011","011101000100","011101000100","011101000100","011100110100","011101000101","100101111000","100001111001","100001111001"),
		("100110001010","100110001010","100110001010","100001100111","100001010100","100001000011","011101000011","100001000100","100001010100","100001000011","011000110011","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","011101000100","011101000101","100001010110","011101010101"),
		("100110001010","100101111000","100101100101","011101000011","011101000011","100001000100","011101000011","011101000011","011101000011","011000110010","010100100010","010000100010","010000100001","010000100001","010000100001","010000100001","010000100001","010000100010","010100100010","010100100010","010000100010","010000100001","010000100001","011000110011","011000110011","011000110011","011000110011"),
		("100101110111","100101100101","011101000011","010100100010","010100100010","010100100010","010000100001","010000100010","010000100001","010000100001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100001","001100100001","010000100001","010000100010","010000100001","001100100001","001100100001","010000100001","010100100010","011000110011","010100100010","010000100010"),
		("100001010100","011101000011","010100100010","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100001","010000100010","010000100010","010000100001","001100100001","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","010100100010","010100100010","010000100001"),
		("011100110011","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010000100001"),
		("011000110010","010100100010","010000100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100010","010000100010","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010000100010","010000100001"),
		("010100100010","010100100010","010000100001","010000100001","010000100001","001100100001","001100100001","010000100001","001100100001","001100100001","010000100001","010000100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100100001","001100100001","010000100001"),
		("011000110011","010100100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001"),
		("011101000101","011000110011","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("100001010110","011000110011","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("100101111000","011000110011","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100001","010000100010","010000100010","010000100001","010000100001","010000100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001"),
		("100110001010","100001010110","010100100010","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100010","010100100010","010100100010","010100100010","010100100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101010101100","100110001001","011000110100","010000100010","010000100010","010100100010","010100110010","010100110010","010100110010","011000110011","011000110011","011000110100","011000110100","011000110100","011000110011","010100110011","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001","001100010001"),
		("101010011100","101010001010","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011000110100","011000110011","011000110011","010100100010","010100100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001","001100010001"),
		("101010101100","100110001001","100001010101","011101000100","011101000100","011100110100","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011101000100","011100110100","011000110011","010100100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101010011100","100101100111","100001000101","011101000100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000100","011000110011","010100100010","010000100010","010000100010","010000100001","010000100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101100","100101100111","011101000100","011101000100","011101000100","011000110100","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","100001000101","100001000101","011000110100","011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101100","100101100111","011101000100","011101000100","011000110100","011000110011","011000110011","011100110011","011000110011","011100110011","011000110011","011000110100","011101000100","100001000101","100001000101","011100110100","011000110011","010100100010","010000100010","010000100010","010000100010","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101100","100101100110","011101000100","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","011101000100","011000110011","010100110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001"),
		("101010101100","100001010110","011100110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","011101000100","011000110011","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001"),
		("101010101100","100001010101","011000110011","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","011101000101","011000110100","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001"),
		("101010001010","011101000100","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","011101000100","011000110011","010100100010","010000100010","010000100010","010100100010","010100100010","010000100010","010000100010","010000100001","010000100001"),
		("100001101000","011000110011","011000110011","011000110011","011000110011","011000110011","010100110011","010100100010","010100100011","011000110011","011000110011","011000110011","011101000101","100001000101","100001000101","100001000101","011101000101","100001000101","011100110100","010100110010","010100100010","010100100010","010100100011","010100100010","010100100010","010000100010","010000100010"),
		("101010011011","011001000100","011000110011","011000110011","010100100010","010100100010","010100100010","010000100010","010100100010","010100100010","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","011101000101","100001000101","100001000101","011100110100","010100110011","010100110011","010100110011","010100110011","010100110011","010100110011","010100100010"),
		("101110101101","100001101000","010100100010","011000110011","011000110011","010100110011","010100100010","010100100010","010100100010","010100100010","010100110010","011000110011","011000110011","011100110100","100001000101","100001000101","011101000101","100001000110","100001000101","011101000100","011000110011","010100110011","010100110011","010100110011","010100110011","010100110011","010100110011"),
		("101110111101","101110101100","011101000101","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010000100010","010100100010","010100100010","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001000101","011101000101","011000110011","011000110011","011000110011","010100110011","010100110011","010100110011","010100110011"),
		("101110111110","101110101101","100001100110","011000110100","011000110100","011000110100","011000110011","010100110010","010100100010","010100100010","010100100010","010100110010","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001000101","100001000101","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011"),
		("101110111110","101110101100","100001010101","011000110011","011000110100","011000110100","011000110011","011000110011","011000110010","011000110011","011000100010","011000110011","011000110011","011000110011","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","011101000101","011000110100","011000110011","011101000100","011100110100","011000110011","011000110100"),
		("101110111110","100101111001","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001000101","100001000101","100001010110","100001010110","011100110100","011100110100"),
		("101110101100","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100101010111","100001010110","100001000101","011000110011"),
		("100001100111","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","100001010101","100001000110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","011000110011"),
		("011100110100","011101000100","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","011101010101","011101000100"),
		("100001010110","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001000101","011101000100","011100110100","011101000101"),
		("101110101100","100001010110","011000110011","011000110010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","011101000100","011101000101","100001010110","100001010110","100001010110","100001010111","100001010110","100001010110","011101000100","011000110011","011000110011","011101000100"),
		("101110101101","100110001001","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011000110011","011000110011","011000110011","011100110100","011100110100","011101000100","011101000100","100001010110","100001010110","100001010110","100001010111","100001010110","100001010110","011000110011","011000110011","011000110011","011100110100"),
		("101110111110","101010101100","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","010000100010","010000110011","010100110100","010101000100","010101000100","011001000100","100001100111","100001100111","100001010110","100001010110","100001010111","100001010111","100001010110","011000110100","011101000100","011101000101","100001000101"),
		("101110111101","101110101101","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010000110011","001100110011","010000110100","010101000100","010101000100","010101010101","011101100111","011101010110","100001000110","100001010110","100001010111","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110101101","100101101000","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","010101000100","010000110011","010000110011","001100110011","001100100011","010101000100","011001010101","010101000100","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110111101","101110111110","101010011011","011101000100","011000110011","011000110010","010100100010","011000110010","010100100010","011000110100","010100110100","010000110100","010001000100","010000110011","010000110011","010001000100","011001010101","011001000100","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110"),
		("101110101101","101110111101","101010101100","100001010110","011000110011","011000110011","011000110011","011000110011","011000110011","011001000100","010000110011","010000110011","010000110100","010000110100","010000110011","010101000100","011001010101","011001010101","100001010110","100001010110","100001010110","100001010110","100001000101","100001010110","100001010110","100001010110","100001010110"),
		("101010011100","101010011100","100110011011","100001101000","011000110011","011000110011","011000110011","011000110011","011000110011","011001000100","010000110011","010000110011","010000110011","010000110011","010000110100","010101000100","011001010101","011101010101","100001000101","100001000101","100001010110","100001010110","011101000101","011101000101","100001000101","100001000101","100001010110"),
		("101010011011","101010011011","100110001010","100001111000","011001000100","010100110011","010100110011","010100100010","010100100010","010100110100","010000110011","001100110011","001100110011","001100110011","010000110011","010101000100","011001010101","011001010101","011101000100","011101000100","011101000101","011101000101","011101000100","011000110100","011101000100","011101000100","100001000101"),
		("100110001010","100110001010","100001111000","100001111000","011001000100","010100100011","010100100010","010000100010","010000100010","010000110011","001100100010","001100100010","001100100010","001100100011","001100110011","010000110100","010101000100","010101000100","011000110100","011000110100","011101000100","011001000100","011000110100","011000110011","011000110100","011000110100","011101000100"))
	-- 16
	,

		(	("101010011100","101010101100","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001","100001111001","100110001010","100110001010","100110001010","100010001001","100001111001","100010001001","100110001001","100110001010","100110001010","100110001010","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101110101100","101010101100","101110101100","101010101100","101010101100","101010101100","101010011100","101010011100","100110001010","100001111001","100001111001","100110001010","101010011011","100110011011","100110001010","100110001010","100110001010","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100010001010","100010001010"),
		("101110101100","101010101100","101010101100","101010101100","101010101100","101010011100","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100110001010","101010011011","100110011011","100110011011","100110001010","100110001010","101010011011","101010011011","101010011100","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010"),
		("101110101101","101110101101","101110101100","101110101100","101010101100","101110101100","101010101100","101010101100","101010011100","100110001010","100010001010","100010001010","100110011011","101010011011","101010011011","101010011011","101010011011","101010011011","101010101100","101010101100","101110101100","101110101100","101110101100","101110101100","100110001010","100110001010","100110001010"),
		("101010011100","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110001010","100110001010","100010001010","100010001001","100001111001","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010"),
		("100110001010","100110001010","100110001011","100110011011","100110011011","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100010001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010"),
		("100110001011","100110011011","100110011011","100110011011","100110011011","100110001010","100010001010","100010001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100010001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010"),
		("100110011011","100110011011","100110011011","100110011011","100110001011","100110001010","100010001010","100010001010","100010001001","100001111001","100001111001","100001111001","100010001001","100010001001","100010001001","100001111001","100001111001","100001111001","100010001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010","100110001010"),
		("100110011011","100110011011","100110011011","100110011011","101010011011","101010011011","100110011011","100110011011","100101111001","100001111000","100001100111","100001100111","100001100111","100001100111","011101010110","011101010101","100001010110","100001100111","100101111001","100110001010","100110011010","100110001010","100110011011","100110011011","100110001010","100110001010","100110001010"),
		("100110011011","100110011011","100110011011","100110001011","100110001011","100110011010","100110001001","100001100110","100001000100","011101000011","011100110011","011100110011","011100110011","011000110011","010100100010","010100100010","011000110010","011000110011","011101000100","011101000101","100001100111","100110001010","100110001010","100110001010","100010001001","100010001010","100110001010"),
		("100110011011","100110011011","100110001010","100110001001","100101111000","100101100110","100101010101","011100110011","011000110011","011000110010","010100110010","011000110011","011000110011","011000110010","010100100010","010100100010","010100100010","010100100010","011000110011","011000110011","011101000100","100001010110","100001100110","100001100111","100001100111","100001111000","100110001010"),
		("100110001011","100110001010","100101111001","100101100110","100101100101","100101100101","011101000011","010100100010","011000110011","011100110011","011101000011","011101000011","011101000011","011000110011","010100100010","010100100010","010100100010","010100100010","010100100010","011000110010","010100110010","011000110011","011100110100","011100110100","011000110011","100001010101","100101111001"),
		("100110001010","100101111000","100101010101","100101010100","100101010100","011100110011","010100100010","001100100001","010000100001","010000100001","010000100001","010000100001","010100100010","010100100010","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010100100010","010100100010","010100100010","011000110011","011101000101","100001100110"),
		("100110001001","100101100101","011101000011","011000110011","011000110010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010000100010","010000100010","010100100010","010100100010","010000100010","011000110011","011101000100"),
		("100101111000","100001010101","011100110011","010100100010","010100100010","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","010000100001","010000100010","010000100010","001100100001","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100001","010000100010","011000110100"),
		("100001010101","011000110011","010100100010","010100100010","010100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100010","010000100010","010100100010","010100100011","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","001100100001","001100100001","001100100001","010100100010"),
		("100001100111","010100110011","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010000100001","010000100010","010000100010","010000100001","010000100010","010000100001","001100100001","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100010001","001100100001"),
		("101010011011","011101000101","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001"),
		("100110011010","100001010110","011000110010","010100100010","010000100010","010000100001","001100100001","001100100001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001"),
		("101010011011","100001010110","011000110011","010100100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101010011011","100101111000","011000110011","010100100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101101","101010011011","100001010110","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010000100010","010000100010","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101101","101110101100","100101111001","011000110100","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000100010","010100100010","010100110011","010100110011","010100100011","010100100010","010000100010","010000100010","010000100010","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001"),
		("101110101101","101010101100","100101111000","011101000100","011000110011","010100110011","010100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000100","011101000100","011100110100","011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001","001100010001","001100010001"),
		("101110101101","101010001010","100001010101","011101000100","011000110100","011000110011","011000110011","011000110011","011000110100","011000110011","011101000100","011101000101","011101000101","100001000101","100001000101","100001000101","100001010101","011101000100","011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100010001","001100010001"),
		("101110101101","100101111000","011101000100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","100001000101","100001000101","100001000101","100001010110","100001000101","011000110100","010100110011","010000100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001"),
		("101010101100","100001100111","011100110100","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001000101","100001000101","100001010110","100001000101","011100110100","010100110011","010100100010","010100100010","010000100010","010000100001","001100100001","001100100001","001100100001"),
		("101010101100","100001100111","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","100001000101","100001000101","100001000101","100001010110","100001000101","011000110100","010100100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001"),
		("101010101100","100101100111","011101000100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","100001000101","100001000101","100001000101","100001010110","100001000101","011000110011","010100110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100010001","001100010001"),
		("101010011011","100001010110","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001000101","100001000101","100001010110","100001000101","011000110100","010100110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100010001"),
		("100110001001","100001010101","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011000110011","011000110011","011000110100","011101000101","100001000101","100001010110","100001000101","011000110100","011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001"),
		("100001010101","011101000100","011000110011","011000110011","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110100","011000110100","011000110011","011100110100","100001000101","100001000101","100001010110","100001000101","011000110100","010100110011","010100100010","010000100010","010000100010","010000100001","010000100001","001100100001","001100100001"),
		("011001000100","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000101","100001000101","100001000101","100001010110","100001010110","011101000100","010100110011","010000100010","010000100010","010000100010","010000100010","010000100010","010000100001","010000100001"),
		("100101111000","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010000100010","010100100010","010100100010","011000110011","011100110100","011101000101","100001000101","100001000101","100001000101","100001010110","100001010110","100001000101","011000110011","010000100010","010000100010","010100100010","010100100010","010000100010","010000100010","010000100010"),
		("101010011011","011001000100","010100100010","011000110011","011000110011","011000110011","010100100010","010000100010","010000100010","010000100010","010100100010","011000110011","011000110100","011101000101","100001000101","100001000101","100001010110","100001010110","100001010110","011101000101","011000110011","010100100010","010100100011","010100110011","010100100010","010100100010","010100100010"),
		("101010011011","011101010101","010100100010","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","011000110011","010100110011","010100100010","010100100010","011000110011","011101000101","100001000101","100001000101","100001010110","100001010110","100001010110","011101000100","010100110011","010100110011","010100110011","010100110011","010100110011","010100110011"),
		("101010001010","100001010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","010000100010","010000100010","010100100010","010100100010","010100100010","011000110011","011100110100","100001000101","100001000101","100001010110","100001010110","100001010110","011101000101","011000110011","010100110011","010100110011","010100110011","011001000100","010100110011"),
		("100101110111","100001010101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010000100010","010000100010","010100100010","010100110011","011000110011","011000110011","011101000101","100001010110","100001010110","100001010110","100001010110","100001000101","011000110011","010100110011","010100110011","010100110011","010100110011","011000110011"),
		("100001010110","100001010101","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011100110100","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","011000110100","010100110011","010100110011","010100110011","011000110011","011000110011"),
		("100101100110","011101000101","011100110100","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","011101000100","011000110011","011000110100","011000110100","011000110011","011100110100"),
		("100001010101","011101000100","100001010110","100001010110","100001000101","011000110011","011000110011","011000110011","011101000100","010100110011","010000100010","010100110011","010101000100","011001000100","011001000100","011101010101","100001100111","100001010110","100001010110","100001010110","100001010111","100001010110","011101000101","100001010110","100001000101","011000110011","011100110100"),
		("011100110100","011101000101","100001010110","100001010110","100001010110","011100110100","011000110011","011000110011","011000110100","010000110011","010000110011","010000110011","010001000100","010101000100","010101000100","011001100110","011101100111","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100101010111","100001010110","011101000100","011000110011"),
		("011000110100","011000110100","011000110011","011100110100","100001000101","011000110100","011000110011","011000110011","011000110011","011001000100","010101000100","010000110011","010000110011","001100110011","010000110011","011001010110","010101000100","011101010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","011101000100","011000110011"),
		("011100110100","011000110100","010100110010","010100100010","011000110011","011000110011","010100100010","010100100010","011000110011","011000110100","010000110011","010000110100","010000110100","010000110011","010000110011","011001010101","010101000100","011101010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","011101000100","011100110100"),
		("011101000101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100110100","010000110011","010000110100","010000110100","010000110011","010000110011","011001010101","011001010101","011101010110","100001000110","100001010110","100001010110","100001010110","100001000101","100001000101","011101000100","011101000100","100001010110"),
		("100001010101","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100110100","010000110011","010000110011","010000110011","010000110011","010101000100","011001010101","011001010101","100001010110","100001000101","100001000101","100001010110","100001010110","011101000101","011000110100","011000110011","011101000100","100001010110"),
		("011101000101","011000110011","011000110011","011000110011","011000110011","010100110011","010100100011","010000100010","010100110011","010100110011","001100110011","001100110011","001100110011","010000110011","010000110011","011001010101","011001010101","011101010101","011101000101","011101000100","011101000101","011101000101","011000110100","010100100010","011000110011","011000110011","011101000101"),
		("011001000101","010100100010","010100100010","010100100010","010000100010","010000100010","010000100001","010000100001","010000100010","010000110011","001100100010","001100100010","001100100010","001100110011","010000110011","010101000100","010101000101","011001000100","011000110100","011000110100","011101000100","011101000100","010100110011","010100100010","011000110011","011000110100","011101000100"))
	-- 17
	,

		(	("101010011100","101010101100","101010011011","101010011011","101010011011","101010011011","101010011011","100110011011","100110011011","100110001010","100001111001","100001111001","100001111001","100110001010","100110001010","100110001010","100010001001","100001111001","100010001001","100110001001","100110001010","100110001010","100110001010","100110011011","100110001010","100001111001","100001111001"),
		("101110101100","101110101100","101010101100","101110101100","101010101100","101010101100","101010101100","101010101100","101010101100","100110001010","100001111001","100001111001","100110001010","101010011011","100110001011","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100010001010","100010001010"),
		("101110101100","101010101100","101010101100","101010101100","101010101100","101010101100","101010011011","101010001010","100101111001","100101100110","100101100101","100001010110","100101110111","100101111000","100101111000","100110001001","100110001010","100110001010","101010011011","101010011011","101010011100","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010"),
		("101110101101","101110101101","101110101100","101110101101","101010011011","100110001001","100001010110","100001010101","011101000100","011100110011","011101000011","100001010100","100001000100","100001000011","100001010100","100101100101","100101100110","100101100111","100101111000","100110001001","101010011011","101010101100","101110101100","101110101100","100110001010","100110001010","100110001010"),
		("101010011100","101010011100","101010011011","101010001010","100101100110","011101000011","010100100010","011000110010","011000110011","011100110011","100001000011","100001000011","011000110011","011100110011","100001000011","011101000011","011101000011","100001000100","100001010101","100101100110","100101110111","100110001010","101010011011","101010011011","100110001010","100110001010","100110001010"),
		("100110001010","100110001010","100101111000","100101100101","100001010100","011000110010","010100100010","100001000100","100001000011","100001000011","100001000011","011000110011","011000110011","011000110011","010100100010","010000100001","010000100001","011000110011","011000110011","011101000100","100001010101","100101100110","100101111000","100010001001","100110001010","100110001010","100110001010"),
		("100110001011","100101111001","100101010101","100101010100","100001000100","011000110010","100001000100","100101010100","011100110011","011000110010","011000110010","010100100010","010000100010","010000100001","010000100001","001100100001","001100100001","010000100010","010100100010","010100100010","011101000100","100001010110","100101100111","100001100111","100001100111","100110001001","100110001010"),
		("100110001010","100101100110","100001000011","100001000100","011101000011","011101000011","100001000011","011101000011","010100100010","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010100110011","011000110011","011000110011","011000110100","011101000100","011101010110","100001111000"),
		("100101100110","011101000011","011000110011","010100100010","010100110010","010100100010","010000100010","010000100001","010000100001","001100100001","001100100001","001100100001","001100010001","001100010001","001100010001","001100010001","001100010001","001100010001","001100100001","001100100001","010000100001","010100100010","011000110011","011101000100","011000110011","010100110010","100001010101"),
		("100101100101","011000110010","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100100010","011000110011","011101000101","011101000101","010100110011","010100110011","011101000101"),
		("100001010100","011000110010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","010000100010","010000100010","010000100010","010100110011","011000110011","011101000100","011101000100","011101000100","011000110011","011000110011","011101000101"),
		("011000110011","010100110010","010000100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","010000100010","010100100010","010100100010","010100100010","010000100010","010000100010","010100100010","010100110010","010100100010","010100100010","011000110011","011000110011","011000110100","011000110011"),
		("011000110010","010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100110011","011000110011","011000110011","011000110011"),
		("010100100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100100010","010100110011","010100110011","010100110011"),
		("010100100010","010000100001","010000100001","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100100010","010000100010","010000100010","010100100010"),
		("011000110011","010100100010","010100100010","010000100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100010","010100100010","010000100010","010000100001","010000100010"),
		("011000110011","010100100010","010000100010","010000100010","010000100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100010","010100100010","010100100010","010100100010","010000100010","010000100010"),
		("011000110011","010100100010","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","001100100001","001100100001","001100100001","001100100001","001100100001","001100100001","010000100001","010000100001","001100100001","010000100001","010000100010","010100100010","010100110011","011000110011","011000110011","011000110011","010100110011","010000100010","010000100010"),
		("010100100010","010100100010","010100100010","010100100010","010100110011","010100110011","010100110011","010100110011","010100110011","010100110010","010100100010","010000100010","010000100010","010000100010","010100100010","010100110011","011000110011","011101000100","011101000101","011101000101","100001010110","100001010110","100001010110","100001010101","011000110100","010100100010","010000100010"),
		("010100100010","010100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001010110","100001010110","100101100111","100101100111","100101100111","100101100111","100101100111","100101100111","011101000101","010100110011","010100100010"),
		("010100100010","010100110011","011000110011","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011101000100","011101000101","100001010110","100001010110","100001010110","100001010111","100101100111","100101101000","100101101000","100101100111","100101100111","100101100111","100001010110","011000110011","010100110011"),
		("010100100010","011000110011","011000110011","011000110011","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011000110100","011101000100","011101000100","011101000101","100001010101","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101100111","100101100111","100101100111","100001010110","011000110100","010100110011"),
		("010100100010","011000110011","011000110100","011000110100","011000110011","011000110100","011000110100","011000110011","011000110100","011000110100","011101000100","011101000100","011101000100","011101000100","011101000101","100001000101","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101100111","100101100111","100001010110","011000110100","010100110011"),
		("010100110011","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000100","011101000100","011101000100","011101000100","011101000101","011101000101","100001000101","100001010101","100001010110","100101010111","100101010111","100101100111","100101100111","100101010111","100001010110","011000110100","011000110011"),
		("010100110011","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110100","011000110011","011101000100","011101000100","011101000101","100001000101","100001000101","100001000101","100001000101","100001000101","100001010110","100101010111","100101010111","100101010111","100101100111","100101010111","100001010110","011101000100","011000110011"),
		("011000110011","011000110011","011000110100","011000110100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000101","011101000101","100001000101","100001000101","100001000101","100001010110","100001010110","100001010111","100101010111","100101010111","100101010111","100101010111","100101010111","100001010110","011000110100","011000110011"),
		("011000110011","011000110011","011000110011","011000110011","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011101000100","100001000101","011101000100","011101000101","100001000101","100001010110","100001010110","100101010111","100101010111","100101010111","100101010111","100101010111","100101010111","100001010110","011000110100","011000110011"),
		("011000110100","011000110100","011000110100","011000110011","010100110011","010100110011","010100110011","010100110011","010100110011","011000110011","011000110100","011101000100","011101000101","011101000100","011101000100","100001000101","100001010110","100001010110","100101010111","100101010111","100101010111","100101010111","100101010111","100101010111","100001010110","011000110100","011000110011"),
		("011101000100","011101000100","011000110011","010100110011","010100100010","010100100010","010000100010","010000100010","010000100010","010100100010","010100110011","011000110011","011000110100","011000110011","011000110011","011100110100","011101000101","100001000101","100001010110","100001010110","100101010110","100101010111","100101010111","100101010111","100101010111","011101000100","011000110011"),
		("011101000101","011101000100","011000110100","011000110011","011000110011","011000110011","010100110011","011000110011","010100100010","010100100010","010100100010","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011101000101","100001010110","100001010110","100101010111","100101010111","011101000100","011000110100"),
		("100001010101","011101000100","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100100010","010100100010","011000110011","011000110011","011101000100","011000110011","011000100011","011000110010","010100110010","011000110011","011000110011","011000110100","011101000100","100001010110","100101010111","100101100111","011101000100","011101000100"),
		("100101100101","011101000100","011000110011","011000110011","011000110011","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011000110011","100001000101","100001010110","011101000101","011000110011","011000110011","011000110011","011000110100","011101000101","100001000101","100001000101","100001010110","100101100111","100101101000","011101000101","100001010110"),
		("100001010101","011101000100","011000110011","011000110011","011000110011","010100100010","010100110010","010100100010","011000110011","011000110011","011000110011","011000110011","100001010110","100101010111","100101010110","011101000101","011000110011","011000110011","011000110100","011101000101","100001010110","100001010110","100101010111","100101101000","100101111000","100001010101","100101100111"),
		("100001010101","011000110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011100110100","100001010110","100101100111","100101100111","100001010110","011101000101","011101000100","011101000101","100001010101","100101010111","100101100111","100101100111","100101111000","100101111000","100001010101","100001000101"),
		("011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110","100101100111","100101100111","100101100111","100001010110","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101111000","100101111000","100001010110","011101000101"),
		("011101000100","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100101100111","100101100111","100101100111","100101100111","100001010110","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101111000","100101111000","100001010111","100001010110"),
		("100001000101","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000101","100101010111","100101100111","100101100111","100001010110","100001010110","100001010110","100001010110","100001010110","100001010110","100101100111","100101100111","100101100111","100101100111","100001100111","100101111000"),
		("100001010110","011100110100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","100001000101","100101100111","100101100111","100101010111","100001010110","100001000110","100001010110","100001010110","100001010110","100001010110","100101010111","100101100111","100101100111","100101100111","100101111000","100110001010"),
		("100101111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","100001010110","100001010110","100001010110","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100001010111","100101100111","100101100111","100101100111","100110001001","101010011011"),
		("100101111000","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","011000110100","011101000100","100001000101","100001000101","100001010110","100001010110","100001010110","100001010110","100001010110","100101100111","100101111001","100110001010","100110001010","101010011011"),
		("100110001001","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011101000100","011000110011","010000100010","010100110011","010100110100","010101000100","010101000100","011001010101","100101111000","100001010110","100001010110","100001010110","100001010110","100001010111","100101111000","100110001010","101010011011","101010011011","101010101100"),
		("101010001010","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010100110011","010000110011","010000110011","010000110100","010001000100","010101000100","011001010110","011101100111","100001010110","100001000110","100001010110","100001010110","100101010111","100101111000","100110011011","101010101100","101010011100","101010101100"),
		("101010011010","011101000101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011001000100","010101000100","010000110011","010000110011","001100110011","001100100011","011001010101","010101000101","011101010110","100001010110","100001010110","100001010110","100101100111","100101111000","101010011011","101010101100","101010101100","101110101101"),
		("101010011011","100001010110","011000110011","011000110011","011000110011","011000110010","010100100010","010100100010","011000110011","011001000100","010000110011","010001000100","010000110100","010000110011","010000110011","010101010101","010101000101","011101010110","100001010110","100001010110","100001010110","100101100111","100110001001","101010011011","101010011100","101010101100","101110101100"),
		("100110001001","100001010101","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110100","010000110011","010000110100","010000110011","010000110100","010000110011","011001010101","011001010101","100001010110","100001000110","100001010110","100001010110","100101101000","100001111001","101010011011","101010011100","101010011100","101110101100"),
		("011101010101","011101000100","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","010101000100","010000110011","010000110011","010000110011","010000110011","010000110100","011001010101","011001010101","100001010110","100001000101","100001000101","100001010110","100001111000","100001111001","101010011011","101010011011","101010011011","101110101100"),
		("011101000101","011101000100","011000110011","011000110011","011000110011","010100110011","010100100011","010100100010","010100110010","010100110100","001100110011","001100110011","001100110011","010000110011","010000110011","010101010101","011001010101","011101010110","011101000101","100001000101","100001010110","100001100111","100001111001","100110001010","100110001011","100110011011","101010011011"),
		("011000110100","010100110011","010100100010","010100100010","010000100010","010000100010","010000100010","010000100010","010000100010","010000110011","001100100010","001100100010","001100100010","001100100011","010000110011","010101000100","010101000100","011001010101","011101000100","011101010101","011101010101","011101010110","100001100111","100001111001","100001111001","100001111001","100010001001"))
	-- 18
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010011011","101010011100","101010011100","101010011100","101010101100","101010011011","100110001010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001010","100110011011","101010101100","101010101100","101010101100","101010101100","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110011010","100110001010","100101110111","100101110111","100101111000","100101111000","100110001001","101010011010","100110001010","100110001010","100110001010","100110001010","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001010","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011011","100101100111","100001000011","011100110011","011000110010","011000100010","011000110010","011101000101","100101111000","101010011011","101010101100","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010001010","100001000100","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","100001010101","101010011011","101010101100","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","101010001010","100101100110","011100110011","010100100010","010100100010","010100100010","010100100010","010100110011","011000110011","011000110011","100110001001","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","101010011011","101010001001","100001010100","011000110011","011101000100","011101000101","100001010101","100001010110","100101100110","100001010110","011000110011","100101111000","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100110001010","101010011100","101010011010","011101000011","011101000100","100001010101","100001010101","100101100110","100101100110","100101100110","100101100110","011101000100","100001100111","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100110001010","100110001010","101010001010","011101000100","011101000100","011101000101","011101000100","100001010101","100101100110","100101010110","100101100110","011101000101","100001111000","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","100010001001","100110001010","011101010101","011101000100","011101000100","011101000100","011101000100","100001010101","011101000101","100001010101","100001010110","100001111000","100110011011","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011010","101010011011","100001111001","100001111000","100001010110","011101000100","011101000100","011101000100","011101000100","100001010110","100101010110","100101010110","100101100110","100001111000","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100010001010","100110001010","100101111001","100001000101","011101000101","011101000101","011101000100","011101000100","100001010101","100101100110","100101100110","100101100110","100110001001","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","100001100110","011101000101","011101000100","011101000100","011101000100","100001010101","100101100110","100101100110","100101100111","100110001001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011100","101010011011","100110001010","100110001010","101010011011","101010011011","100110011011","100001111001","100001100111","011101000101","011101000100","011101000100","100001010101","100101010110","100101100110","100001111000","100001111001","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011011","100110011011","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100110001010","100001010101","011101000100","011101000101","100001010110","100101100110","100101100110","100001111000","100110001010","100110001010","100001111001","100110001010","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100110001010","101010011010","100001100110","100001010110","011101000101","100001010101","100001010110","100001010110","100001100111","011101100111","101010011010","100110001001","100001111001","100110001010","100001111001","100001111000","100001111000"),
		("100010001001","100110001010","101010011100","101010011100","100110011011","100110001010","100110001010","100010001001","100001111001","100001111001","100110001010","100110001010","011101010101","011001010101","011101000101","011101000101","100001010110","100001010110","100001100111","010000110011","010101000100","011101100110","100001100111","100001111000","100001111001","100001111001","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110011011","100110001010","100110001010","100110001001","100001111001","100110001001","101010011010","100110001001","011001010101","011001010101","011101010101","100001000101","100001010110","100001100111","011101100111","001100100010","001100100010","001100100010","010000100010","010101000100","011001010101","011101100111","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110011011","100110001010","100010001010","100110001010","100001111001","100001111001","100110001010","100101111000","011001010101","011001010101","011101010101","100001000101","100001010101","100001100111","011101100110","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","010000110011"),
		("101010011011","100110001010","100110001010","101010011011","100110011010","100010001001","100010001001","100110001010","100010001001","100001111000","011101100111","011101010101","011001010101","011001010101","011101000101","011101000100","011101000101","100101111001","011101100111","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010"),
		("101010101100","100110001010","100110001010","101010011011","100110001010","100010001001","100001111001","100010001001","100101111001","011101010101","010000100010","010100110011","011101010110","011001010101","011101000101","011101000100","100001100111","100001111001","010000110100","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110011010","100110001010","100110011010","100110001010","100110001010","100001111001","100010001001","100001111000","011001000100","010000100010","001100100001","010000110011","100001100111","011101100111","100001010110","100001010110","100001111000","011001010110","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001010","100110001010","100110001001","100010001001","100001111000","100001100110","011000110100","001100100001","001100100001","001000100001","001100100010","100001100111","011101100111","011001010101","011001010101","011001000101","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001010","101010011011","100110001010","100001111001","100001111001","011101010110","010000100010","001100100010","001000100010","001000100010","001000100010","001000100001","011101010110","011101100111","010101000101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","101010011011","101010011011","100110001001","100101111001","010101000100","001100100001","001000100010","001000100010","001000100001","001000100001","001000100001","010101000101","011001010110","010101000100","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("101010011100","101010011011","101010011011","100110011010","100101111001","010101000100","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010"),
		("101010011011","101010011011","101010011011","101010011010","100001111001","011001000101","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010000110100","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010"),
		("101010101100","101010101100","101010011011","100110001001","100001111001","011101010110","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010000110011","010101000100","010000110100","001100100010","001100100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","101010011100","100110001001","100001111000","100001111001","011101100111","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010000110011","010001000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100010","001000100010"),
		("100110001010","100110001010","100110001001","100110001001","100001111001","011101100111","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","001100110011","010000110100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010"),
		("100110001010","100110001001","101010011010","101010011010","100001111001","011101100111","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","001100110011","010000110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010"),
		("100110001010","100110001010","101010011011","100110011010","100001111001","100001111000","010000110011","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","001100110011","010000110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100010"),
		("100110001010","100110001010","100110011010","100110011010","100001111001","100001111000","011001010101","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","001100100010","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001001","100110001010","100010001001","100001111000","011101100110","001100100010","001000100001","001000100001","001000100001","001000010001","001100110011","001100100010","001100110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000010001","001000100001","001000100010"),
		("101010011011","101010011011","100110001001","100010001001","100010001001","100001111000","011001000100","001000100001","001000010001","001000010001","001000010001","001000010001","001100110011","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","000100010001","001100110010","001000100010"),
		("101010011100","101010011011","100110001010","100110001001","100001111001","100001111000","010000110011","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000010001","001000010001","001000100001","001000100001"),
		("100110001010","100110001010","100110001010","100001111000","100101111000","011101010110","010000100010","001000100001","001000010001","001000010001","001000010001","001000010001","001100110010","001100100010","001100100010","001100100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","000100010001","001000010001","001000010001","001000100001"),
		("100110001010","100110001010","100101111000","100001010110","100001010110","100001010101","010000110011","001100100001","001000010001","001000010001","001000100001","001000100001","001100110010","001100100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000010001","000100010000","001000010001","001000100001","001000100001"),
		("100110001010","100110001001","011101010101","100001000101","100001010110","100001010110","010100110011","001000100001","001000010001","000100010001","001000100001","001000010001","001100110011","001100100010","001000100001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100001","001000010001","000100010000","000100010000","001000010001","001000100001","001000100010"),
		("100110011010","100101111001","011101000100","011101000100","100001010101","100001010110","011001000100","001000010001","000100010001","000100010001","001000100001","001000010001","001100110011","010000110011","010000110011","001100100010","001000100001","001000100010","001000100001","010000100011","010000100010","001100100001","001000010001","000100010001","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100001010110","011000110100","011101000101","100001010110","011101000100","001000010001","000100010000","000100010001","001000010001","001000010001","001100110011","010101000100","010101000100","010000110011","001000100001","001000100001","001000100001","010100110011","011100110100","011000110011","010100110011","001000100010","001000100001","001000100010","001000100010"),
		("100110001010","100110001001","100001111000","011101010110","011101000100","011101000100","010000100010","001000010001","001100110011","001000100010","000100010001","001000010001","001100110011","010101000100","010101000100","010000110100","001000100010","001000100001","001000010001","011000110011","011101000100","011101000100","011101000100","010000100011","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100001111001","100001111000","010000110011","001100010001","010000110011","011101100110","011101100111","001000100010","000100010001","001000010001","001100110011","010101000100","010101000100","010101000100","001000100010","001000010001","000100010000","010100110010","011101000101","011101010101","011101000101","010100110100","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","010101000101","001100110011","011101111000","100110001001","011101010110","001100100010","000100010001","000100010001","001100110011","010101000100","010101000100","010101000100","001000100010","000100010001","000100010000","001100100010","011101000100","011101000101","011101000101","011001000100","001000100010","001100100010","001100100010"),
		("011101100111","011101100111","100001100111","100001110111","100001100111","011101100111","100001111000","011101100110","010000110011","001100100010","000100010001","000100010000","001100110010","010100110100","010101000100","010101000100","001100100010","000100010001","000100010000","001000100001","010100110011","011101000100","011101000100","010100110100","001000100010","001000100010","001000100010"),
		("011101100110","011101100110","011101100110","011101100110","011101100110","011101100111","011101100111","010101000100","001100100010","001000100001","000100010001","000100010000","001100100010","010000110011","010000110100","010000110100","001100100010","000100010001","000100010000","000100010000","001100100010","010100110011","010100110011","010000100010","001000100001","001000100001","001000100010"))
	-- 19
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100010001001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","100110001001","100101100110","100101100110","100001100110","100001100110","100001111000","100110001010","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100010001001","100110001010","100110001001","011101000011","011000110010","010100100010","010100100010","010100100010","011000110011","100001100111","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100101111000","100101010101","011000110010","010000100001","010000100001","010000100001","010100100010","010100100010","011000110011","100101111000","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110011011","100110001001","100101010101","011101000011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000100010","011101010110","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001010","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011100","101010011010","100001010100","011000110010","011101000100","011101000101","100001010101","100001010101","100001010110","100001010110","011000110100","011101010110","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011010","011101000100","011000110011","100001010101","100001010101","100001010110","100101100110","100101100110","100101100110","100001000101","011101010110","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011100","101010011010","011101000100","011100110100","011101000101","011101000100","100001010101","100101100110","100101100110","100101100110","100001010101","011101010110","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010101100","101010011011","011101010101","011101000100","011101000100","011101000100","011101000100","100001010101","011101000101","011101000101","100001010101","100110001001","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100110001010","101010011011","101010011011","101010101100","100110001001","100001010101","011101000101","011101000101","100001010101","011101000100","100001010101","100101010110","100001010110","100001100110","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010101100","100101111000","100001000100","100001000101","011101000101","011101000101","011101000100","100001010101","100101100110","100101100111","100101100111","101010011010","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","100010001001","100110001010","101010011011","100110001001","100001010110","011101000101","011101000100","011101000100","011101000100","100001010101","100101100110","100101100110","100101111000","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011010","101010011011","100001111001","100001111001","100010001001","100001111001","100110001001","100001100111","011101000100","011101000100","011101000100","100001010110","100101010110","100101100111","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100010001010","100110001010","101010011010","100110001010","100010001001","100110001010","100001100111","011101000100","011101000101","100001010101","100101100110","100101100110","100001111000","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011011","100010001001","100110001001","100001010110","011101000100","011101000100","011101000100","100001010110","100101010110","100001101000","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011100","101010011011","100110001010","100110001010","101010011011","101010011011","100110011011","100010001001","100001111000","100001111000","100001010110","011101000100","011101000100","011101000100","100001010110","100001010110","011101010110","011001010110","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011011","100110011011","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100110001010","100101111000","100001010101","011101000101","011101000100","100001010101","100101100110","100101010111","011101010110","001100100011","010101000100","100001111000","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100110001010","100110001010","100110001010","100001111001","100001111000","100001100111","100101100111","100001010110","011101010101","011101000100","100001010101","100001010110","100001100111","011001010101","001100100010","001100100010","001100100010","010100110100","011101010110","100001111000","100001111001"),
		("100010001001","100110001010","101010011100","101010011100","100110011011","100110001010","100110001010","100010001001","100001111000","011101010110","010100110011","010100110011","011101010110","011001010101","011101010101","011101000101","011101000100","011101010101","100101111000","010101000100","001100100010","001100100010","001000100010","001000100001","001000100001","001100100010","010101000100"),
		("100010001010","100001111001","100110011011","101010011011","100110011011","100110001010","100101111001","011101010110","010100110011","010000100010","001100100001","010000110011","011001010101","011001010101","011101010101","011101000100","011101010101","100001111000","100110001001","010000110100","001100100010","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001"),
		("100110011011","100010001001","100110001010","101010011011","100110001010","011101100111","011001000100","010000100010","001100100010","001000100010","001000100001","001100100010","011001010101","011001010101","011101100110","100001010110","100101111000","100110001001","011001010101","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","100110001010","100110001010","101010011011","100110001001","010000110011","001100100010","001100100010","001000100010","001000100010","001000100010","001100100010","011001010101","011001010101","011001010110","011001010101","011001010110","011001010110","001100110011","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010"),
		("101010101100","100110001010","100110001010","101010011011","100001111001","010000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","011001010101","011001010101","010101000101","010101000101","010101000100","001100100010","011001000100","011001000100","010100110011","001100100010","001000100010","001000100010","001000100010","001000100010"),
		("100110011010","100110001010","100110011010","100110001010","100001111000","001100100010","001000100010","001000100010","001000100001","001000100001","001100100001","001100100001","010000110011","011101100110","010101000101","011001000101","010101000101","010000110011","010000110011","100001010101","100001000101","011101000101","011001000100","001100100010","001000100010","001000100010","001000100010"),
		("100110001010","100110001010","100110001010","100110001001","100001111000","001100100010","001000100010","001000100001","001100100001","001100100001","001000100001","001000100001","010000110011","100001100111","011001010101","010101000100","010101000100","001100110011","010101000100","100001010101","011101000101","011101010101","011101000100","001100100010","001000100010","001000100010","001000100010"),
		("100110001010","101010011011","100110001010","100010001001","011101100111","001100100010","001000100001","001100100010","001000100010","001000100010","001000100010","001000100001","010101000100","100001111000","011001010101","010101000100","010000110011","001100100010","011001000100","100001000101","100001000101","100001010101","011101000100","001000100010","001000100010","001000100010","001000100010"),
		("101010011011","101010011011","101010011011","100110001001","011101100111","001100100010","001100100001","001000100010","001000100010","001000100001","001000100001","001000100001","010000110011","011101100110","010101000101","010001000100","010000110011","001100100010","010000100010","011100110100","011101000101","100001010101","011101000100","001100100010","001000100010","001000100010","001000100010"),
		("101010011100","101010011011","101010011011","100110011010","011101100111","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010101000100","010001000100","010000110011","001000100010","001000100010","010100110011","011101000100","100001010101","011101000100","001100100010","001000100010","001000100010","001000100010"),
		("101010011011","101010011011","101010011011","101010011011","011101100111","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010001000100","010000110100","001100110011","001000100010","001000100010","001100100010","011000110011","011101000101","011101000100","001100100010","001000100001","001000100010","001000100010"),
		("101010101100","101010101100","101010011011","100110001001","100001111000","001100100010","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110100","010000110100","001100100010","001100100010","001100100010","001000100010","001100100010","010100110011","010100110011","001100100010","001000100001","001000100010","001000100010"),
		("101010011011","101010011100","100110001001","100001111000","100001111000","010000100010","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010001000100","010000110011","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","001000100010","010000110011","001000100010","001000100010"),
		("100110001010","100110001010","100110001001","100110001001","100001111000","010000110011","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110011","010000110011","001100100010","001000100010","001000100010","001000100010","001000010001","001000100001","001000100001","001000100010","011001010101","001100100010","001000100001"),
		("100110001010","100110001001","101010011010","101010011010","011101100111","001100100010","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110011","001100110011","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000010001","001000010001","001000100010","001000100010","001000100010"),
		("100110001010","100110001010","101010011011","101010011010","011101010110","010000100010","011001000100","010000100010","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110011","001100100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110011010","100110011010","011101010110","100001010101","100001010101","011000110011","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010000110011","001100110010","001000100010","001000100001","001000010001","001000010001","000100010001","001000010001","000100010000","000100010000","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001001","100110001010","100001111000","100001010101","100001010101","011101000100","001100100010","001000100001","001000100001","001000010001","001100100010","010000110100","010000110011","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","001000010001","001000100001","001000100010"),
		("101010011011","101010011011","100110001001","100010001001","100001010110","011100110100","100001010101","100001000101","010000100010","001000010001","001000010001","001000010001","001100100010","010000110011","001100100010","001100100010","001000100001","001000010001","001000010001","000100010001","000100010000","001000100001","001100100010","001000010001","000100010001","001100110011","001000100001"),
		("101010011100","101010011011","100110001010","100110001001","100001100111","011101000100","011101000101","100001010101","010000100010","000100010001","001000010001","001000010001","001100110011","010000110011","001100100010","001100100010","001000100001","001000100001","000100010001","000100010000","000100010000","001000100001","001100110011","001000010001","001000010001","001000100001","001000100001"),
		("100110001010","100110001010","100110001010","100110001001","100001100111","011000110100","011101000100","011101000100","010000100010","001000100001","001000010001","001000010001","001100110010","010000110011","001000100010","001000100001","001000100001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001"),
		("100110001010","100110001010","100110001010","100110001001","100001111000","011001000100","010000100010","010000110010","011101100111","010000110011","001000010001","001000010001","001100110010","010000110100","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001010","100110001001","100110001001","011101100111","010000110011","011101100110","100101111000","001100110011","001000100001","001000100001","010000110011","010101000100","010101000100","001100100010","001000100001","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","000100010000","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001010","100110001001","100001111001","100001111001","100001111001","100110001001","100001110111","001100100010","001000100010","001000100010","010101000100","010101000101","010101000100","001100100010","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100010"),
		("100110001010","100110001010","100110001001","100110001001","100001111000","100001111000","100001111000","100110001001","011101010110","001100110011","001100110011","001100100010","010101000100","010101000101","010101000100","001100110011","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100001111001","100001111000","100001111000","100001111000","100110001001","011001010101","001100100010","010000110011","001100110011","011001010101","010101000101","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100001111001","100001111000","100001111000","100001111000","100001111000","100101111001","010101000101","001100100010","001100100011","010000110011","010101010101","010101000101","010101000100","010000110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","100001110111","100001111000","100001111000","100001111001","010000110100","001000100010","001100100010","010000110100","010101000101","010101000101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","001000100010"),
		("011101100111","011101100111","100001100111","100001110111","100001110111","100001111000","100001111000","011101100111","001100110011","001000100010","010000110011","010101000100","010101000100","010101000100","010101000101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("011101100110","011101100110","011101100110","011101100110","011101100110","011101100111","011101100111","011001010110","001100100010","001000100010","010000110011","010000110100","010000110100","010001000100","010101000100","010000110100","010000110011","001100100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100001","001000100001","001000100010"))
	-- 20
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100001111001","100001111001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011010","101010001010","101010001010","101010011010","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010001010","100101100110","100001010100","100001000100","011101000100","011101010101","100001100111","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001001","100101100110","011000110010","010100100010","010100100010","010100100010","010100100010","011000110011","100001100111","100110001001","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110011010","100110001010","100101100110","100001000100","010100100010","010000100001","010000100001","010000100001","010000100001","010100100010","011000110011","100001111000","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011100","101010001010","100101010101","011100110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000110011","011000100010","100001100111","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011010","011101000100","011100110011","100001010101","100001010101","100001010110","100101100110","100101100110","100101010110","011000110011","100001100111","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010101100","101010001001","011000110011","011101000100","011101000101","100001010101","100001010110","100101100110","100101100110","100101100110","011101000100","100001100111","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010101100","101010001010","011100110100","011101000100","011101000100","011101000100","100001010101","100001010110","100001010110","100101010110","011101000100","100101111000","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100110001010","101010011011","101010011011","101010101100","100110001001","100001010101","100001000101","011101000100","011101000100","011101000100","100001010110","011101000101","100001010101","100001010110","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100110001010","100110001010","101010011011","101010011011","100001010110","100001010101","100001010101","011101000101","011101000101","011101000100","100101100110","100101100110","100101010110","100101100111","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","100010001001","100110001010","101010011011","100101100111","100001000100","011101000101","011101000100","011101000100","011101000100","100001010110","100101100110","100101100110","100101100111","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011010","101010011011","100001111001","100001111001","100010001001","100001111001","100001100111","100001010101","011101000100","011101000100","100001010101","100101010110","100101100110","100101100111","100001111000","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100010001010","100110001010","101010011010","100110001010","100010001001","100110001001","100001010101","011101000100","011101000100","100001000101","100101010110","100101100110","100101111000","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010011011","100010001001","100001111000","011101000101","011101000100","011101000100","100001010110","100101100110","100101100111","100101111001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","100110011011","100010001001","100001111001","100001100111","011101000100","011101000100","011101000100","011101000101","100001010110","100001100111","100001111001","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100110001010","100110001010","101010011011","101010011011","100110001010","100010001001","100110001001","100001100111","011101000100","011101000101","011101000101","100001010101","100101010110","100001100111","100110001001","100110001010","100001111000","100110001001","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100010001001","100110001010","100110001001","100001111000","100001100111","100101111000","100001100110","100001010101","011101000101","011101000101","100001010110","100001010110","100001100111","011001010101","100110001001","100110001001","100001111001","100110001010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010101100","100110011011","100110001001","100101111000","011101100111","011001000100","010100110011","010100110011","100001100110","011101010101","011001010101","011101000101","011101000101","100001010101","100001010110","100001111000","010000110011","010000110011","011001010101","100001100111","100101111001","100010001001","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100001100111","011101010101","010100110011","010000100010","001100100010","001100100010","010000100010","100001010110","011001010101","011001010101","100001010110","011101000100","011101000101","100001111000","011101100111","001100100010","001100100010","001100100010","001100100010","010101000100","011101100111","100001111000","100001111001"),
		("100110011011","100010001001","100110001010","011101100111","010000100010","001100100010","001100100001","001100100001","001100100010","001000100010","001100100010","100001100110","011001010101","011001010101","100001010110","011101000101","100001100111","100110001001","011101100111","001100100010","001100100010","001000100010","001000100010","001000100001","001000100010","010000110011","011101100111"),
		("101010011011","100110001010","100001111001","010101000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","011001000101","011001000101","011001010101","011101010110","100001111000","100110001001","100001111001","010000110100","001100100010","001100100010","001000100010","001000100010","001100100010","001100100010","001000100001","001100100010"),
		("101010101100","100110011010","100001111000","010000100010","001000100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001100110010","010101000100","011001010101","011001010101","011001010101","100001111000","011001010101","001100100010","001100100010","001000100010","001000100001","001100100010","011101000100","011101010101","010101000100","001100100010"),
		("100110011010","100110001010","100001100111","001100100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001","001100100001","001100100010","011001010101","011001010110","011001000101","011001010101","011001010101","010000110011","001000100010","001000100010","001000100010","001000100001","001100110011","100001010101","100001010110","100001010110","011001000100"),
		("100110001010","100001111001","011001000101","001100100010","001000100010","001100100010","001000100010","001000100001","001100100001","001100100001","001000100001","001100100010","011101100110","011101100110","010101000101","011001010101","010101000101","001100110011","001000100010","001000100010","001000100010","001000100001","010000110011","011101000101","100001010110","100001010110","011001000100"),
		("100110001010","100001111000","001100100010","001000100001","001000100001","001000100001","001100100001","001100100010","001000100010","001000100010","001000100010","001000100010","011101100111","011101100110","010101000101","010101000101","010101000100","001100100010","001000100010","001000100001","001000100001","001000100001","001100100010","011000110100","100001010101","100001010110","010100110011"),
		("101010011011","011101100111","001000100001","001000100001","001000100001","001000100001","001100100001","001000100010","001000100010","001000100001","001000100001","001000100001","011001010101","011001010101","010101000100","010101000101","010000110100","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","010100110011","100001000101","100001010101","010000110010"),
		("101010011011","011101100110","001000100001","001000100001","001000100001","001000100001","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","010000110011","010101000101","010101000100","010101000100","010000110011","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","010000110011","011101000101","100001010101","010000100010"),
		("101010011011","011001010101","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","001100100010","011101000100","100001000101","010000110011"),
		("100001111000","010101000100","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","001000100001","010000110011","010101000100","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","001000100001","001100100010","010000110011","001100100010"),
		("010101000100","001100100010","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","010100110011","011101000100","011001000100","011001000100","010101000100","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100100010","001100100010"),
		("001100100010","001100100001","001000100001","001000100001","001000010001","001000100001","001100100001","001000100001","010000110011","011101000100","011101000101","011101000100","011001000100","010000110011","010000110100","010000110011","001100100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001"),
		("001100100001","010000100010","001100100010","001100100001","001100100001","010000110011","001100100001","001100100001","011000110011","011101000100","011101000101","011101000101","011001000100","010000110011","010000110011","010000110011","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001"),
		("001100100001","001100100010","001000100001","001000100001","001100100010","001100100010","001000100001","001100100001","011000110011","011101000100","011101000100","011101000100","010100110100","010000110100","010000110011","001100110011","001000100010","001000100001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","001000010001","001000010001","000100010001"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000100010","010100110011","010000100010","001100100010","010000110011","010001000100","010000110011","001100100010","001000100010","001000100001","001000010001","001000010001","000100010001","001000010001","000100010000","000100010000","001000010001","001000010001","000100010000"),
		("001100100001","001000100001","001000100001","001000100001","001000100001","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001100110011","010000110100","010000110011","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","000100010001","001000010001","001000010001","000100010000"),
		("010101000101","001100100010","001000100001","001000100001","001000100001","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010000110100","010000110011","001100100010","001000100001","001000010001","001000010001","000100010001","000100010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010000"),
		("101010011011","100110001010","011101100111","011001010101","011001010101","011001010110","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010000110011","010000110011","001100100010","001000100001","001000100001","000100010001","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000010001","001000010001"),
		("100110001010","100110011010","100110001010","100110001001","100101111000","100001100111","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001"),
		("100110001010","100110001010","100110001010","100110001001","100001111000","100001100111","001100100010","001000100001","001000010001","001000100001","001000100001","001000100001","001100110011","001100110011","001100100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001"),
		("100110001010","100110001010","100110001010","100110001001","100001111000","100001111000","010000110011","001000100001","001000100001","001000100001","001000100001","001000010001","001100110011","001100100010","001000010001","001000010001","001000100001","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","000100010000","001000010001","001000010001","010101000100"),
		("100110001010","100110001010","100110001010","100110001001","100001111001","100001111000","001100110011","001000100001","001000100001","001000100001","001000100001","001000010001","001100110011","001100110011","001100100010","001000100010","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001100110011"),
		("100110001010","100110001010","100110001001","100110001001","100001111001","100001111000","001100110010","001000100001","001000100001","001000100001","001000010001","001000010001","001100110011","010101000100","010101000100","010000110011","001000100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010"),
		("100110001010","100110001001","100010001001","100001111001","100001111001","100001111000","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100110011","010001000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010"),
		("100110001001","100010001001","100001111001","100001111000","100001111000","100001111000","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100110011","010000110100","010101000101","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100010"),
		("100001111000","100001111000","100001111000","100001111000","100001111000","011101100111","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100110010","010000110011","010101000101","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010"),
		("011101100111","011101100111","100001100111","100001110111","100001111000","100001100111","001100110011","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","001100100010","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","001000100001"),
		("011101100110","011101100110","011101100110","011101100110","011101100110","011101100110","001100110011","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","001100100010","010000110100","010000110100","001100100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001"))
	-- 21
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100101111000","101010001001","100110001001","101010011010","101010011011","101010101100","101010011011","100110001010","100110001001","100110001001","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110001001","100101100101","100001000100","011101000011","011000110010","011000110011","100001010110","100110001001","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","100101111000","011000110010","010100100010","010100100010","010100100010","010100100010","010100100010","011101000100","100101111000","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010001001","100001010101","010100110010","010000100001","010000100001","010000100001","010000100010","010100100010","010100100010","011101010110","101010011011","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","100101111000","100001010100","011000110011","011000110100","011101000100","011101000100","100001010101","011101010101","011000110011","011001000101","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","101010011011","100101110111","011101000011","100001010101","100001010101","100101100110","100101100110","100101100110","100101100111","011101000101","011001000100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100110001010","101010101100","100001100111","011000110011","100001000101","011101000101","100001010101","100101100110","100101100110","100101100110","100001010101","011101000100","101010011010","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100110001010","100110001010","100101111001","011101000100","011101000100","011101000100","011101000100","100001010101","011101000101","100001010110","100001010101","011101010110","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100110011011","100010001001","100101111000","100001010101","011101000100","011101000100","011101000100","100001010110","100001010101","100001010110","100001010110","100001100111","100001111001","100110011010","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011010","101010011011","100001111001","100001010110","100101100110","100001000101","011101000100","011101000100","100001010110","100101100110","100101100110","100101100110","100101100111","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100010001010","100110001010","100101111000","100001010101","100001010101","011101000101","011101000100","100001010101","100101100110","100101100110","100101010110","100101111000","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100110001010","101010011011","101010011011","100101111001","100001010101","011101000101","011101000101","100001010110","100101100110","100101100110","100101111000","100110001010","100110001001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","100110011011","100110001001","100001010110","011101000101","011101000100","100001010110","100101100110","100101100110","100110001001","100010001001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100110001010","100110001010","101010011011","101010011011","100110001010","100001111001","100001010101","011101000100","011101000101","100001010110","100101010110","100001100110","100001111000","100001111000","100110001010","100110001010","100001111000","100110001001","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100001111001","100110001001","100110001010","100001111000","100101111000","100001010110","100001010101","011101010101","100001000101","100001010110","100001010110","100001111000","100110001001","101010011011","101010011011","100110001001","100001111001","100110001010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011100","100110001010","100010001001","100010001001","100001111001","100001111000","100001111000","100101100111","011101010101","011001010101","011001010101","100001010110","100001010110","100001010110","100001100111","100001111000","101010011011","101010011011","100110001010","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110001010","100110001001","100001111001","100001100111","011101010110","011101010101","100001100111","011101010110","011001010101","011001010101","100001010110","100001010110","100001010110","011101100110","010000110011","011001100110","100110001001","100110001010","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110001001","100001100111","011101000101","010100110011","001100100010","010000100010","100101111000","100001100111","010101000101","011001010101","100001010101","100001010101","100001100111","011001010110","001100100010","001100100010","001100100010","010001000100","011101100110","100101111000","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100001111000","100001100111","011001000100","010000110010","001100100010","001000100010","001000100001","001100100010","100101111000","100001100111","010101000101","011001010101","011101000101","011101010110","100110001001","011001010110","001100100010","001100100010","001100100010","001000100010","001000100010","010000110011","011001010110","100001111000","100001111001"),
		("101010011100","100001111001","010100110100","010000100010","001000100010","001100100010","001000100010","001000100010","001000100001","010000110011","100101111000","100001100111","011001010101","011001010101","100001100110","100101111001","100110001010","010101000101","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","010000110011","011101100111"),
		("100110011010","011101010110","001100100010","001100100010","001000100010","001100100010","001000100010","001000100010","001000100001","001100100010","011001000100","011001010110","011101100110","011101100110","100001110111","100110001001","011101100111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010000110011"),
		("100010001001","011001000101","001000100010","001100100010","001000100010","001100100010","001000100010","001000100001","001100100001","001100100001","001100100001","010101000100","100001100111","011001010110","011001000101","011101010110","010000110100","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010"),
		("100110001001","010101000100","001000100010","001000100001","001000100001","001000100001","001100100001","001100100010","001000100010","001000100010","001000100010","010101000100","100001110111","011001010110","011001010101","010101000101","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001100100010"),
		("100110001001","010000110011","001000100001","001000100001","001000100001","001000100001","001100100001","001000100010","001000100010","001000100001","001000100001","010101000100","011101100110","011001010101","011001010101","010101000100","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010","001100100010"),
		("100110001001","001100100010","001000100001","001000100001","001000100001","001000100001","001100100010","001000100010","001000100001","001000100001","001000100001","010000110011","010101000101","011001010101","010101000101","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010"),
		("100001111001","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","011001000101","011001000101","010101000100","010000110011","001000100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100010"),
		("100001111000","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000101","010101000101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001100100010","011000110100","010101000100","001100100010","001000100001","001000100010","001000100010"),
		("100001111000","001100100010","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","011101000100","100001010110","011101010101","010000110011","001000100010","001000100010"),
		("100001100111","001100100010","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000010001","001100100010","010101000100","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","010000100010","100001000101","100001010110","100001010110","011001000100","001000100010","001000100010"),
		("100001100111","001100100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100010","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","010000110011","100001010101","100001010110","100001010110","010100110011","001000100010","001000100010"),
		("011001010101","001100100010","001000100001","001000100001","001000100001","001100100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","010000110011","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","001100100010","011101000100","100001010101","011101000100","001100100010","001000100001","001100100010"),
		("001100100010","001000100001","001000100001","001100100010","011001000100","011001000100","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010000110100","001100110011","001000100001","001000100010","001000100001","001000100001","000100010001","001000100001","011000110011","011101000100","010100110011","001000100001","001000100001","001000100010"),
		("010000110011","001100100010","011001000100","100001010110","100001010110","011000110011","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000100010","011000110011","010100110011","001000100001","001000100001","001000100010"),
		("010000110100","010100110011","011101000101","011101000100","011101000100","011000110100","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","000100010001","000100010000","000100010001","001000100001","001000100001","001000010001","001000100001","001000100010"),
		("010000110011","010100110011","011100110100","011000110011","011101000100","011000110100","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000100001","000100010001","000100010000","000100010000","000100010001","001000100001","001000010001","001000100010","001000100010","001000100001"),
		("001100100010","010000100010","011000110011","011100110011","011101000100","011000110100","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000100001","001100100010","001000100010"),
		("010101000100","001100100010","010000100010","011000110011","011000110011","001100100010","001000010001","001000100001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000010001","001000100001","001000100010"),
		("100110001001","011001010101","001100100010","010000100010","001100100010","000100010001","001000010001","001000100001","001000010001","001000010001","001000100001","001000010001","010000110011","001100110011","001000100010","001000100001","001000100001","001000100010","001000010001","000100010001","001000010001","001000010001","001000100001","000100010000","000100010001","001000010001","001100110011"),
		("100110001001","100110001001","011001010101","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","001100100010","001000100001","001000010001","001000100001","001000100010","001000100001","001000010001","001000100001","001000010001","010101000100","011001010101","010001000100","011001010101","100001111000"),
		("100110001010","100110001010","100001111000","001100100010","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","001000010001","010000110011","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","001000010001","010101000100","100110001001","100110001001","100110001001","100110001001"),
		("100110001010","100110001001","011101100111","001000100001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","010000110100","010101010101","010101000100","001100100010","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","010000110011","100101111000","100110001001","100110001001","100110001001"),
		("100110001001","100010001001","011001010110","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","010000110100","011001010101","010101000101","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100100010","011101100111","100110001001","100110001001","100110001001"),
		("100001111000","100001111000","011001010101","001000100001","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000110011","011001010101","010101000101","010000110011","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","010101000100","100001111001","100001111001","100001111001"),
		("011101100111","100001100111","010101000101","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","011001010101","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010001000100","100001111000","100001111000","100001111000"),
		("011101100110","011101100110","010000110100","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010101000100","010101000100","010000110011","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","010000110011","011101100111","011101100111","011101100111"))
	-- 22
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110001010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110011010","100110011011","100010001010","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010001010","101010001010","101010001001","100101111000","100110001001","100110011010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","100101111000","100101100101","100001010100","011100110011","011000110011","011101000100","100101100111","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001001","100001000100","011000110011","011000110010","010100100010","010100100010","011000110011","011000110011","100001010101","100110001001","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100101111000","011100110011","010000100001","010000100001","010100100010","010000100001","010100100010","010100100010","010100100010","100001100111","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100101110111","011101000011","011000110011","011000110011","011001000100","011101000100","100001010101","011101000100","010100100010","011101010101","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100101100111","100101010101","100001010101","100001010110","100101100110","100101100110","100101100110","100001010110","010100110011","011101010101","100110001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100101100111","100101010110","100001010101","100001010101","100001010110","100101100110","100101100110","100101010110","011000110011","011101010101","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110011011","100110001001","100001010110","011101000100","011101000100","100001010101","011101000101","100001010101","100101010110","011100110100","100001010110","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100101111001","100001010101","011101000100","011101000100","100001010110","100001010101","100001010101","100001010110","011101000100","100001111000","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100101111000","100001010110","011101000101","011101000101","100001010110","100101100110","100101100110","100101100110","100001010110","100101100111","101010011011","100110001010","100110001001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100110001010","100110001010","100110001001","100001010110","011101000100","011101000100","100001010110","100101100110","100101100110","100101100110","100101100110","100101111000","100110011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100110001010","100110001010","101010011010","100101110111","011101000100","011101000100","100001010101","100101010110","100101100110","100101100110","100101111000","100110001010","100110001001","100001111000","100110001010","100110001010","100001111000","100110001010","101010011010","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100010001001","100110001010","100101111001","011101000100","011101000100","100001010101","100001010110","100101100110","100101100110","100101111000","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100001111001","100110001010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011100","100110001010","100010001001","100010001001","100001111001","100001111000","100001010101","011101000100","011101010101","011101010101","011001010101","100001100110","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110001010","100001111001","100001111001","100101111001","100001111000","011101010101","011101000100","011101000101","011001010101","011001010101","100001100110","100001111000","100110001001","101010011010","100110011010","101010011011","101010011011","101010001010","100101111001","100001111000","100001111000","100001111000","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110001010","100001111001","100001111001","100110001001","100101111000","011101000100","011100110100","011101010101","011001010101","011001010101","100001010110","100001100111","011001010101","100001111000","100110001001","101010011011","101010011011","101010011010","100101111001","100101111001","100010001001","100001111000","100001111000"),
		("101010011011","100010001001","100001111001","101010011010","100110001010","100001111001","100001111000","011101010110","011101010110","011101000100","011101000100","011101000101","011001010101","011001010101","100001010110","100001100111","010000110011","001100100011","010000110100","011001010110","100001111000","100001111000","100001111001","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100001111001","100110001010","100110001001","100001010110","010100110011","001100100010","011001000100","100001100111","011101000100","011101000101","011001010101","011001010101","011101010110","100001111000","010000110011","001100100010","001100100010","001000100010","001000100010","001100110010","010101000101","100001100111","100110001001","100001111000","100001111000"),
		("100110001010","100010001001","100110001010","100001111000","011101000101","010000100010","001000100001","001000100001","010000110011","100101111000","100001100110","011101010101","011101100110","011101010101","100001100111","100110001001","010001000100","001100100010","001100100010","001000100010","001000100010","001000100001","001000100001","001000100010","010101000100","100001111000","100001111000"),
		("100001111001","100001111000","011101010110","010100110011","001100100010","001000100010","001000100010","001000100001","010000110010","100001110111","100110001001","100001100111","100001100111","100001100111","100110001001","100001111001","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100001111001"),
		("011101100111","010100110100","001100100010","001000100001","001000100001","001000100001","001100100001","001100100010","001100100010","011101100110","011101100111","011101100111","100001111000","100001100111","100001111001","011001010110","001100100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","011001010101","100001111001"),
		("010101000100","001100100010","001000100001","001000100001","001000100001","001000100001","001100100001","001000100010","001000100010","001100100010","010000110100","010101000100","011101010110","011001010101","010101000101","001100110011","001000100010","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","010101000100","100101111001"),
		("010000110011","001100100010","001000100001","001000100001","001000100001","001000100001","001100100010","001000100010","001000100001","001000100001","010000110011","011001010101","011001000101","011001010101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010001000100","100110001001"),
		("010000110011","001100100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100110010","010101000100","011001000101","010101000101","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","100101111001"),
		("010000100010","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","011001000101","010101000100","010000110100","010000110011","010100110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100001111000"),
		("001100100010","001100100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010101000100","010101000100","010101000100","010000110011","010000110011","011101000101","100001010110","011001000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000"),
		("001100100010","001100100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","010000110011","010101000100","010101000100","001100110011","010000110011","100001010101","100001010101","100001010110","010100110011","001000100001","001000100010","001000100010","001000100001","001000100010","001100100010","100001111000"),
		("010000110011","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001100110011","010101000100","010101000100","001100110011","010000110011","100001000101","100001010101","100001010101","010100110011","001000100010","001000100001","001000100001","001000100001","001000100001","001100100010","100001111000"),
		("010000110011","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001100100010","010101000100","010001000100","001100110011","010000100010","011101000100","011101000101","100001010101","010100110011","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","100001110111"),
		("010000110011","001100100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000010001","001100100010","010101000100","010101000100","001100110011","001000100001","001100100010","011101000100","011101010101","010100110011","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010101000100"),
		("100001010110","011101000100","001100100010","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","010001000100","010000110100","001100110011","001000100001","001000010001","010100110011","011101000100","010000110011","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010"),
		("100001010110","100001010101","011001000100","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110011","001100110011","001000100001","001000010001","001000010001","001100100001","001000100001","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010"),
		("100001010101","100001010110","100001010110","010000110010","000100010001","001000010001","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110100","010000110011","001000100001","001000010001","001000010001","000100010000","001000010001","001100100010","001000100010","001000100001","001000100001","001000100010","001000100001","001000100001"),
		("100001010101","100001010110","100001010110","011000110100","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","010000110011","010000110011","001100110011","001000100010","001000100001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001000100001"),
		("011101000101","100001010110","100001010110","011001000100","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110011","010000110011","001100110011","001100100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","001100100010"),
		("011000110100","100001000101","100001010101","010000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","010000110011","010000110011","001100110011","001000100010","001000100001","001000100010","001000010001","000100010001","001000010001","001000010001","000100010001","000100010001","000100010001","001000100001","011001010110"),
		("010100110011","010000100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","010000110011","010000110011","001100100010","001000100010","001000100001","001000100010","001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001100100010","011001010110","100110001001"),
		("010000110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","010000110011","001100110011","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100001","010000110100","100001111000","100001100111","100001111000","100110001001","100110001001"),
		("011001010110","001100110011","010000110011","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001100110011","001100100010","001000100010","001000100001","001000100010","001000100001","001000100010","001000100010","001000100001","010000110011","100101111000","100110001001","100110001001","100110001001","100110001001"),
		("100001111001","100001111000","010101000101","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","010000110011","010101000100","010000110011","001100100010","001100100010","001000100010","001000100010","001000100010","001000100001","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001"),
		("100001111000","011101100111","001100100010","001000010001","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000110011","011001010110","011001010110","010101000101","010000110100","001100100010","001000100010","001000100001","001000100010","001000100010","011101100110","100110001001","100001111001","100001111001","100001111001"),
		("011101100111","011001010101","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010000110011","011001010101","011001010101","010101000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100001","010101010101","100001111000","100001111000","100001111000","100001111000"),
		("011101100110","010101000100","001000010001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100110011","010101000101","010101000100","010101000100","010000110011","001100110011","001000100010","001000100010","001000100010","001000010001","010001000100","011101100111","011101100111","011101100111","011101100111"))
	-- 23
	,

		(	("101010011011","101010011011","101010011011","100110011011","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110001010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","101010011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010011011","101010101100","101010101100","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001010","101010011011","101010001001","101010001001","101010001001","101010001010","101010101100","101010011011","100110001010","100110001001","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001010","100110001010","100101100110","100101010101","100001000100","011000110011","011101000011","100001100110","101010001010","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011011","100110011011","100110001010","100101111000","011101000011","010100100010","010100100010","010100100010","010100100010","011000100010","011000110011","100001100111","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110011011","100110001010","100101110111","011100110011","010000100001","010000100001","010000100001","010000100001","010100100010","010100100010","011000110011","100101111000","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110011011","100110011011","100101111000","100001010101","011101000100","011000110011","011001000100","011001000100","011000110011","010100100010","010100100010","011101010110","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101100","100110011011","100110001010","100101111000","100001010101","100001010101","100001010110","100101100110","100101100110","100101100110","011000110011","010000100010","011101010110","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110011011","100110001010","100101100111","011101000101","100001010101","100001010110","100101100110","100101100110","100101100110","011000110011","010100100010","100001100111","101010011011","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100110011011","100110001010","100001010110","011101000100","011101000101","011101000101","100001010101","100101100110","100101100110","011000110011","010100110011","100101111000","101010011011","100110001010","100110001001","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100110001011","100110001010","100001010110","011101000100","100001010101","100001010101","011101000100","100001010110","100101100110","011000110011","011001000100","101010001010","100110011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100110001010","100110001001","100001010101","100001000101","100101010110","100101100110","100001010110","100101100110","100101100110","011101000100","100001100111","101010011010","100110001001","100001111000","100110001010","100110001010","100001111000","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","101010011011","100110001010","100001111001","100001010101","011101000100","100001010101","100001010110","100001010110","100001100110","100101100111","100001010110","100001100111","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100001111001","100110001010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011100","100110001010","100010001001","100101111001","100001010101","011101000100","100001010101","100001010110","100001010110","011001010101","011001010101","100001100110","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111000","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110001010","100001111001","100001111001","100001010110","011101000100","011101000101","100001010101","100001010101","011001010101","011001010101","100110001001","100110001001","100110001001","101010011010","100110011010","101010011011","101010011011","101010011010","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110001010","100001111001","100001111001","100001100111","011101000100","100001000101","100001010101","100001010101","011001000101","011101010110","100110001001","100001111001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011010","100101111001","100101111001","100010001001","100001111000","100001111000"),
		("101010011011","100010001001","100001111001","101010011011","100110001010","100001111001","100001111000","100001010101","011100110100","011100110100","011101000100","011101010101","010101000101","011001010101","100001111000","100001111000","100001111000","100001111000","100110001010","101010011011","101010011011","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001010","100010001001","100110001001","100101111000","011101010110","100001010110","011101000100","011100110011","011100110100","100001010101","100001010110","011001010101","011101100110","100001111000","100001111001","100001111001","100001111000","100001111001","100110001010","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("100110001010","100001111000","011101010110","010100110011","010000110010","010000100010","011101010110","011101010101","011100110100","011101000100","011101000101","100001010110","011101100110","100001100111","010101000101","011101100111","100110001001","100110001001","100001111001","100001111000","100001111000","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("011101010110","010100110011","001100100010","001100100001","001000100001","001000100010","011101010101","100001111000","011101000101","011101000100","011101000101","100001010110","100001100111","100001111000","010000110011","001100100010","010000110011","011101010110","100001111000","100001111001","100110001001","100001111001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001100100010","001000100010","001000100010","001000100001","001000100001","001100100010","100001100111","100110001001","100001100111","100001000101","100001000101","011101000101","100001111000","011101100111","001100100011","001100100010","001000100010","001000100010","001100110011","011001010101","100001111000","100110001001","100010001001","100001111001","100001111001","100001111001","100001111000"),
		("001000100001","001100100010","001000100001","001000100001","001000100001","001000100010","011101010110","100001111000","100001111000","100001100110","011101010110","100001111000","100001111000","011001010101","001100100010","001100100010","001100100010","001100100010","001000100001","001000010001","001100100010","011001010110","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001100100010","001000100001","001000100001","001000100001","001000100001","001100100010","010000110011","010101000100","011001010110","100001100111","100110001001","011101100111","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000010001","011101100110","100110001001","100001111001","100001111000","100001111000"),
		("001000100010","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000101","010101000100","010101000100","011001010110","011001010110","001100100011","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","001000010001","010001000100","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","011001000101","011001010101","011001010101","011001010101","010101000101","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001100100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010101000100","011001010101","011001010101","011001010101","010101000100","001100110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100100010","100001111000","100010001001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110100","011001010101","011001010101","011001010101","010101000100","001100100011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100100010","100001111000","100110001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001100100001","001000100001","001000010001","001100100010","011001000100","011101000101","011101010101","011001010101","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001100100010","100001111000","100110001001","100110001001","100001111001"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010100110011","011101000101","100001010101","100001010101","011101010101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100001","001100110010","100001111000","100110001001","100010001001","100101111001"),
		("001000100001","001000100001","001000100001","001000100001","001000010001","001100100010","011000110100","011101000101","100001000101","100001000101","011001000101","010001000100","010101000100","001100100010","001000100010","001000100001","001000100001","001000100010","001000100010","001000100010","001000100010","001000010001","001100110011","100001111001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000100001","001000100001","000100010001","010000100010","011000110100","011101000100","011101000101","011101000100","010101000100","010000110100","010101000100","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100001","010000110011","100110001001","100110001001","100110001001","100110001001"),
		("001000010001","001000010001","001000010001","001000010001","000100010001","010000100010","011100110100","011000110011","010000100010","010000110011","010001000100","010000110100","010000110100","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100010","001000100001","010000110011","100110001001","100110001001","100001111000","100001100111"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","010000100010","010100100010","001100100001","000100010001","001000100001","010000110011","010101000100","010101000100","001100100011","001000100001","001000100001","001000100001","001000010001","000100010001","001000010001","001000100001","001000100010","001100100010","011101100111","100001110111","011001000100","011101000100"),
		("001000010001","001000010001","001000010001","001100100010","001000100010","001000100001","001000100001","001000010001","001000010001","001000100001","010000110011","010000110011","010001000100","001100110011","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","010000110011","011101000101","011000110011","011101000100"),
		("001000010001","001000010001","001000100001","001100100010","001000100001","001000010001","001000010001","001000100001","001000010001","001000100001","001100110011","010000110011","010000110100","001100110010","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000100010","011000110011","011000110100","011101010101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000100001","001100110011","010000110011","010001000100","010000110011","001000100001","001000010001","001000100001","001000100010","001000010001","000100010001","001000010001","001000010001","001000010001","010100100010","011000110011","011000110011","100001010101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","010000110011","010000110100","001100110011","001000100001","001000010001","001000100001","001000100010","001000100001","001000010001","001000100001","001000010001","001000010001","010100100010","011000110011","011000110011","011101000101"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100010","010000110011","010000110011","001100110011","001000100001","001000010001","001000100001","001000100001","001000010001","000100010001","000100010001","000100010001","000100010000","001100100001","010000100010","010000100010","010100110011"),
		("010101000100","010101010101","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000100001","001000010001","001000100001","010000110011","010000110011","001100100011","001000100010","001000100001","001000100001","001000100001","001000010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010001","001000010001","001000100001"),
		("100001111001","011101100111","001000100010","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001100100010","010000110011","001100100010","001100100010","001100100010","001000100001","001000010001","000100010001","000100010000","000100010000","000100010000","000100010000","000100010000","000100010000","001000100001","010101000100"),
		("100001111000","011101100111","001000100010","001000100001","001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","010000110011","001100110011","010000110011","010000110011","001000100010","001000100001","001000100001","000100010001","001000100001","001100110010","001100110010","001100110010","010001000100","011001100110","100001111000"),
		("011101100111","011101010110","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100100010","010001000100","010101000101","011001010101","010101000100","001100100010","001000100001","001000100001","000100010001","001000100001","011001010110","100001110111","100001111000","100001111000","100001111000","100001111000"),
		("011101100110","011001010101","001000100001","001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","001100100010","010101000100","010101000101","010101000101","010101000100","010000110011","001000100001","001000010001","000100010001","000100010001","001100100010","011001010110","011101100111","011101100111","011101100111","011101100111"))
	-- 24
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101110101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100110001010","100010001001","100010001001","100110001010","100110011011","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001010","100010001010","100010001001","100010001001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110011011","100110001010","100110011011","100110001010","100110001010","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101110101100","100110011011","100110001011","100110001010","100110001010","101010011011","101010011011","101010011011","100110011010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101110101100","100110011011","100110001010","100110001010","101010011011","101010001010","101010011010","101010011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","101010011011","101010101100","100110011011","100110001010","100110001001","100101100110","100101010101","100001010101","100001010101","100101110111","101010011011","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","101010011011","100110011011","100110001010","100110001001","100001010101","011000110011","011000110011","011000100010","010100100010","011000100010","011101000100","100101111000","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101110101101","101010011100","100110011011","100101110111","100001000100","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","100101111000","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101110111101","101110101100","100110001011","100101100111","100001000100","010100110011","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","100001100111","101010011010","100001111001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101110101101","101110111101","101110101101","100110001010","100001010101","100001010101","100001010101","100001010101","100001010101","100001010110","100101010110","011101000101","010100100010","100001100111","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110111101","101110101100","101110101100","101110111110","101110101101","100110001001","100001010101","100001010101","100001010101","100001010101","100001010110","100101100110","100101100110","100101010110","011000110011","100001111000","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110111101","101010101100","100110001010","100101100110","100001010101","011101000100","100001010101","100001010101","100001010110","100101100110","100001010110","011000110011","100110001001","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011100","101110101101","101010101100","100101111001","100101100111","100001000101","011101000100","011101000100","100001010101","011101000100","100001010101","100001010110","011101010101","101010011010","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100101111000","100101100110","100001010101","011101000100","100001010101","100101100110","100001010101","100101010110","100001010110","100001010110","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110011011","100101111001","100101100110","100001000101","011101000100","100001000101","100101010110","100101100110","100101100110","100101010110","100001100111","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100110001010","100110001010","101010101100","101110101100","101010011011","100110001010","100101111000","100001000101","011101000100","011101000101","100001010110","100001010110","100001100110","100101100110","100101111000","100010001001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011100","100110001010","100010001001","100101111001","100001010101","011101000100","011101000100","100001010101","100001010110","011001010101","011001010101","100101111001","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100010001010","100001111001","100110011011","101010011011","100110001010","100010001001","100001111000","100001000101","011101000100","011101000101","100001010101","100001010101","011001010101","011001010101","100110001001","100110001001","100110001001","101010011010","100110011010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110011011","100010001001","100110001010","101010011011","100110001010","100001111000","100101100110","011101000100","011101000100","011101000100","100001010101","100001010101","011001010101","011001010101","100110001001","100001111001","100001111001","100110001010","101010011010","101010011011","101010011011","101010011010","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100010001001","101010011010","100101111000","011101010101","100001010110","011101000100","011100110100","011000110011","100001000101","100001010101","010101000101","011001010101","100001111000","100001111000","100001111000","100001111000","100110001010","101010011011","101010011011","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","011101100111","011001000100","010100110011","010000100010","100001010110","011101000100","011100110011","011100110100","100001010101","100001010110","011001010101","011001010101","011001010110","100001111000","100001111001","100001111001","100001111001","100110001010","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("100001100110","010100110100","010000100010","001100100001","001100100001","001100100010","100001100111","100001100110","011100110100","011101000100","100001000101","100001010101","011101100110","011001010110","001100100010","001100110011","011001010101","100001111000","100001111001","100001111001","100001111000","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001100100010","001100100010","001000100010","001100100010","001000100001","001000100010","011101010110","100101111000","011101010101","011101000101","011101000101","011101010101","100001111000","011001010110","001100100010","001100100010","001000100010","001100110011","011001010101","100001111000","100110001001","100110001001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","011101100110","100110001001","100001111001","100001010110","100001010101","100001111000","100110001001","011001010101","001100100010","001100100010","001100100010","001000100010","001000100001","010000110011","011101100110","100001111001","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001100100010","001000100001","001000100001","001000100001","001000100001","010000110100","010101010101","011001010110","011101010110","100001110111","100110001001","100001111000","010101000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100001","001000100010","011101100110","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001100110010","011001010101","010101000101","010101000101","011101100111","011001010110","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000010001","010101000100","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","011001010101","011001010101","011101010110","011001010110","011001010101","001100110011","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100001","010000110011","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010101000100","011001010101","011001010110","011001010110","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110100","011001010101","011001010101","011001010101","010101000100","001100100011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","100101111000","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100001","010000110011","011001010101","010101000101","011001010101","010101000100","001100100011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","100001111001","100110001001","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001100100010","010000100010","001000100001","001000100001","001000100001","001100100010","011001010101","010101000101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001100110011","100001111001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000100001","010100110011","100001010101","011000110011","001000100001","001000100010","001000100010","001100100010","011001010101","010101000100","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100001","001100100010","100001111000","100110001001","100110001001","100010001001","100101111001"),
		("001000100001","011001000100","011101000101","011101000100","011000110011","001100100010","001000100010","001000100010","001000100010","010101000100","010101000100","010000110100","010101000100","001100100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","001100100010","100001111000","100110001001","100110001001","100110001001","100001111001"),
		("001100100010","011000110100","011000110011","011100110100","011001000100","001100100010","001000100010","001000100010","001000100010","010000110011","010101000100","010000110100","010101000100","001100100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001"),
		("001000100001","011000110011","011000110011","011000110100","011000110100","001100100010","001000100010","001000100010","001000100001","001100100010","010101000100","010000110100","010000110100","001100100010","001000100001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100010","010000110011","100001110111","100110001001","100110001001","100101111001","100001111001"),
		("001000100001","010000100010","011000110011","011000110100","010100110011","001000100001","001000100001","001000100001","001000100001","001100100010","010000110100","010101000100","010000110100","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001000100010","010000110011","011000110100","011101100110","100101111001","100110001001","100010001001","100001111000"),
		("001000010001","001100100001","010100110011","011000110011","001100100001","001000010001","001000100001","001000100001","001000100001","001000100010","010000110011","010000110100","010001000100","001100100010","001000100001","001000100001","001000100001","001000010001","001000010001","001100100010","011000110011","011100110100","011101010101","100001111000","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001100100010","001100100010","001000010001","001000010001","001000010001","001000100001","001000010001","001000100001","010000110011","010000110100","010000110100","001100100010","001000010001","001000100001","001000100001","001000010001","001000010001","010000100010","011000110011","011101000100","011101000101","100001100111","100110001001","100110001001","100001111001"),
		("001000010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","010000110011","010000110011","010000110100","001100100010","001000010001","001000010001","001000100001","001000100001","001000010001","010000100010","011000110011","011101000101","100001010110","100001111000","100110001001","100110001001","100001111001"),
		("001100100010","001000100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000010001","001100110011","010000110011","010000110011","001100100010","001000010001","001000010001","001000010001","001000010001","000100010001","010000100010","011000110011","011101000100","100001100111","100101111000","100110001001","100110001001","100001111001"),
		("001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001100100010","010000110011","010000110011","001100100010","001000100001","001000010001","000100010001","000100010000","000100010000","001000010001","010000100010","010100100010","011101010110","100110001001","100110001001","100110001001","100001111001"),
		("001000100001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000100001","001000100010","001100100010","010000110011","010000110011","001000100010","001000010001","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","010101000101","100110001001","100110001001","100110001001","100001111001"),
		("001000100001","000100010000","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100010","001000100010","010000110011","010000110011","001100100010","001000010001","001000010001","001000010001","000100010000","000100010000","000100010000","001100100010","011101100111","100010001001","100110001001","100010001001","100010001001"),
		("001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","001100100010","010001000100","010101000100","010000110011","001100100010","000100010001","000100010000","001000100010","010101000100","010001000100","010101000101","011101100111","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001100100010","011001010110","010101000100","010000110100","001100100010","001000010001","000100010000","001000010001","011001010101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000100010","010101000101","010001000100","010101000100","001100100010","001000010001","000100010000","000100010000","001100100010","011101100110","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 25
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011100","100010001010","100001111001","100001111001","100110001010","100110011011","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100110001010","100010001001","100010001001","100110001011","100110011011","100110011011","100010001001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110011011","100110001010","100110001010","100110001001","100101111000","100101111000","100101111001","100001111001","100110001010","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110011011","101010011011","101010101100","100110001010","100101110111","100101010101","011101000011","100001000100","011101000100","011101000100","100001010110","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010101100","101010101100","100101110111","100101010100","011000110010","010100100010","010100100010","010000100001","010100100010","010100100010","100001100111","100110011010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010101100","101010001001","100001010100","011000110010","010000100001","010000100001","010000100001","010000100001","010000100001","010100100010","100101110111","100110011010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101101","101110101101","101010011100","100110001010","011001000011","010100100010","010000100010","010000100001","010100100010","010100100010","010100110010","010100110011","011101000100","100110001001","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","101010011011","100110001001","010100110010","010000100001","010000100001","010100110011","011101000100","100001010101","100101100110","100101100110","100101100110","100101111000","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","101010011100","101010011011","011000110011","010000100001","010100100010","011001000100","100001010101","100001010110","100101100110","100101100111","100101100111","100101111000","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100001111001","100001111001","100001111001"),
		("101010011011","100110011011","101110101101","101010011011","011000110011","010000100001","010100100010","011101000100","011101000101","100001010101","100001010110","100101100110","100101100110","100001100111","100110001001","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","101010011011","011000110011","010100100010","010100100010","011101000100","011101000101","011101000101","100001010101","100001010101","100101010110","100101100111","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110111101","101110101100","101010101100","101010101100","100001010110","011100110011","011000110011","011101000100","100001010101","100001010101","100001010110","100001010101","100001010110","100101111000","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101101","101110101100","101010101100","101110101101","100101111000","011101000100","011101000100","011101000100","011101000100","100001010101","100001010110","011101000100","100001010101","100101111000","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101110101100","101110101100","101010011011","101110101101","101010011011","100001010110","011101000100","011101000100","011101000100","011101000101","100001010101","100001010101","100001010110","100101111000","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010011011","101010011011","100101111000","011101000101","011101000101","011101000100","011101000101","100001010101","100001010101","100101010110","100101111000","101010011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100110001010","100110011011","101010011011","101010011100","100110001010","100101111001","100001000101","011101000100","011101000100","011101000100","100001010101","100001010110","100101100111","100001111000","100110001001","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100010001010","100110001010","101010101100","101110101100","100110011011","100101111000","100001000101","011101000100","011101000100","011101000100","011101000100","100001010101","100001100111","100001111000","100001111000","100110001001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100010001001","100110001010","101010011011","101010011011","100001100111","011001000100","011101000100","011101000100","011101000100","011101000100","100001000101","100001010110","011001010101","011001010101","011101100110","011101100111","100001111000","100110001010","101010011011","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100010001010","100010001001","100101111001","011101010110","010000100010","010000100010","011101010110","011101000100","011101000100","011101000100","100001010101","100001010101","011001010101","011001010101","010001000100","001100100010","010000110100","011001010110","100001111001","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110001001","011101100111","010100110011","001100100010","001000100001","001100100010","011101100110","011101010101","011101000100","011101000100","100001010101","011101000101","010101010101","011001010101","010001000100","001100100010","001100100010","001100100010","001100100010","011001010110","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("011001000100","010000100010","001000100010","001000100010","001000100010","001000100001","010101000101","100001111000","011101000101","100001010101","100001000101","011001000100","011001000101","011001010101","010000110100","001100100010","001100100010","001100100010","001100100010","001100100010","100001111000","100110001001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001100100010","001100100010","001000100001","010000110011","100001111000","100101111001","100001100110","011101000101","100001100111","011101100110","011001010101","001100110011","001100100010","001100100010","001100100010","001100100010","001100100010","011001010110","100001111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001100100001","001100100001","001000100010","001100110010","100001100111","100110001001","100001111000","011101100111","011101100111","011101100111","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010101000101","100110001001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001100100010","001100100010","001100100010","001100100010","001000100001","001000100010","001000100010","010101000101","011101100110","011001010110","011101100110","011001010101","011101100110","011001010110","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010101000101","100110001001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100010","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","001100100010","010101000101","011001010110","011001100110","010101010101","011101100111","011001010110","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","010101000100","100001111001","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","010101000100","011001010110","011001010110","010101000100","011001010101","010101000101","001100100010","001100100010","001100100010","001100100010","001000100010","001000100001","010001000100","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010000110011","011001010110","011001010101","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","011001010101","010101000101","010101000100","010101000100","001100110011","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000101","010101000101","010001000100","010000110100","010101000100","010000110011","010000110011","001100100010","001000100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000100","010000110011","010000110011","010101000100","011101000100","011101010101","011101000101","001100100010","001000100010","001000100010","001000100010","100001100111","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100010","010000110011","010001000100","010000110011","001100110011","010100110100","011101000100","100001010101","100001010101","010000110011","001000100001","001000100010","001000100001","011001100110","100110001001","100110001001","100010001001","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000010001","001000010001","001000010001","001000100001","001000100010","001000100010","001100110011","010001000100","001100110011","001100110011","010100110100","011101000100","100001010101","100001010101","010000110011","001000100001","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100010","001000100010","001100100010","010000110100","001100100010","001100100010","010000110011","011000110100","011101000101","011101010101","010000100010","001000100001","001000100010","001000100001","001000100001","011101100111","100110001001","100110001001","100010001001","100101111001"),
		("001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","001000100010","001000100010","001100100010","010000110011","001000100010","001100100010","001100100010","001000010001","010100110011","011101000100","001100100010","001000100001","001000100010","001000100001","001100100010","011101100111","100110001001","100110001001","100110001001","100001111001"),
		("000100010001","001000010001","000100010001","000100010001","000100010000","000100010000","000100010001","001000100001","001000100010","001100100010","010000110011","001000100001","001100100010","001100100010","000100010000","001100100010","010000100010","001000100001","001000100001","001000100001","001000100001","011001010110","100110001001","100110001001","100110001001","100110001001","100010001001"),
		("001000010001","000100010001","000100010001","000100010001","000100010001","000100010000","000100010000","001000010001","001000100001","001100100010","010000110011","001000100010","001100110011","001000100010","001000010001","001000100001","001000010001","001000100010","001000100010","001000010001","001100110011","100001111000","100110001001","100110001001","100110001001","100101111001","100001111000"),
		("001000010001","001000100001","010000100010","001100100010","001000010001","001000010001","000100010001","000100010001","001000010001","001000100010","001100110011","001000100010","001100110011","001100100010","000100010001","001000100001","001000100001","001000010001","001000100010","001100100010","011101100110","100110001001","100110001001","100101111001","100110001001","100010001001","100001111000"),
		("001000100001","010000100010","011000110100","011000110011","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","001100100010","001100110011","001100100010","001000010001","001000010001","001000100001","001100110010","011001010110","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("010100110011","011101000100","100001010101","011101000101","001100100010","000100010001","001000010001","001000010001","001000010001","001000100001","001100100010","001000100010","001100110011","001100100010","001000010001","001000010001","010000110011","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("010000100010","011000110011","011101000100","100001010101","010000100010","000100010001","001000010001","000100010001","001000010001","001000010001","001000100001","001000100001","001100110011","001100100010","001000100001","001000010001","001100110011","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100101111001","100110001001","100110001001","100001111001"),
		("001100100001","011000110011","011100110100","100001000101","010000100010","000100010001","001000010001","001000010001","001000010001","001000100001","001100100010","001100100010","001100110011","001100100010","001000100001","001000100001","001000100001","011101100111","100110001001","100110001001","100110001001","100110001001","100110001001","100101111001","100110001001","100110001001","100001111001"),
		("001000010001","001100100001","011000110011","011101000100","001100100010","000100010001","001000010001","000100010001","001000010001","001100110011","010101000101","010000110011","010000110011","001100100010","001000100001","001000100001","001000100001","010101000101","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000100001","000100010001","001000100001","001000100001","001000010001","001000010001","001000010001","000100010001","001000010001","010000110011","011001010101","010101000100","010000110011","001100100010","001000100001","001000100001","001000100001","010000110011","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000100001","000100010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","010000110011","011001010101","010101000100","010000110011","001100100010","001000100010","001000100010","001000100001","001100110011","100001111000","100110001001","100110001001","100110001001","100010001001","100010001001","100110001001","100010001001","100010001001"),
		("001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","010000110011","011001010101","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","011101100111","100010001001","100001111001","100001111001","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("000100010001","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","010001000100","011001010101","010101000101","010000110100","001100100010","001000100001","001000100010","001000100010","001000100001","011001010101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010000","001000100010","001000100001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","010101000100","010101010101","010101000101","010000110011","010000110011","001000100010","001000100001","001000100001","001000010001","010001000100","011101100111","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 26
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100101111000","100101110111","100001100111","100001100111","100001111000","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100101111001","100101100110","100001000100","011000110011","010100100010","010100100010","010100110010","011000110011","100101111000","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110011011","100110001010","100101100101","011101000011","010100100010","010000100001","010000100001","010000100001","010000100010","010100100001","011000110011","101010011010","101010101100","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001011","100110011011","100101100111","011101000011","010100100010","010000100001","010000100010","010000100001","010000100001","010000100001","010000100001","011000110011","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","100110001001","011001000011","010000100001","010000100001","010000100001","010100100010","011000110011","011000110011","011001000100","011000110011","100001100111","100110011010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","100001100111","010100100010","010000100001","010100100010","010000100001","011000110011","100001010101","100101100110","100101100111","100101100111","100101111000","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100001100110","010100100001","010000100001","010000100001","010100100010","011101000100","100001010101","100101100110","100101100111","100101100111","100101111000","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110011010","100001111001","100001111001","100010001001"),
		("101110101101","101010101100","100110001010","011101010101","010000100001","010000100001","010000100001","010100100010","011101000100","100001000101","100001010101","100001010101","100001010110","100101100111","101010011010","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","101010011011","011101010101","010100100001","011000110011","010100100010","010100110011","011101000101","100001010101","100001010101","100001010101","100001010101","100001100111","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101110101100","100001111000","011000110011","100001000101","011101000100","011100110100","011101000101","100001010101","100001010110","100101100110","100001010110","100001100111","100110001001","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","101010011010","011000110011","011101000100","011101000101","011101000100","011101000100","011101000101","100001010101","100101100110","100001010101","100001010110","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110111101","101010101100","101010101100","101010101100","100001100111","011100110011","011101000100","011101000100","011101000100","011101000101","100001010110","100001010110","100001010110","100101111000","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101010101100","101010011100","101010011011","101110101101","100110001001","011101000101","011101000100","011101000100","011101000100","011101000100","100001010101","100001010101","100001010101","100110001001","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011011","101010101100","101010011011","101010011010","100101111000","100001000101","011101000100","011101000100","011101000100","011101000100","011101000101","100001010101","100101100110","100110001001","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("100110001010","101010011011","100101111001","011001000101","100001010101","011101000100","011101000100","011101000101","011101000101","011101000100","011101000101","100001100110","100001100111","100001111000","100110011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100001111001","100001100111","010100110011","001100100001","011101010101","011101000101","011101000100","011101000101","011101000101","100001010101","100001100111","011101100111","100001100111","100001111000","100110001001","101010011011","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("010101000100","001100100010","001000100010","001000100010","011001000101","100001100110","011101000100","100001000101","100001010101","100001010101","100001100111","011001000101","011001010101","011101100111","011101100111","100001111000","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","100110011010","100010001001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","010000110011","100001111000","011101010101","100001000101","100001010110","011101000101","100001111000","011101100111","011001000101","011001010101","010101000100","001100100011","010101000101","100001111000","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100001","010000110010","100001111000","100001111001","100001010110","100001000101","011101000101","100110001001","100001111000","011001000101","011001010101","010101000100","001100100010","001100100010","001100110011","100001111000","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001100100010","001000100010","001100100010","011101100111","100110001010","100001111000","011101010110","100001111000","100110001010","011001010101","010101000101","011001010101","010101000100","001100100010","001100100010","001000100010","011001010110","101010011011","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001000100010","001000100010","010000110011","011001010110","011001010110","011101010110","011001100110","011001010110","010000110011","010101000100","011001010101","010101000100","001100100010","001100100010","001100100010","010101000100","100110001010","101010011010","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001100100010","001000100001","010001000100","011001010110","011001010101","011001010101","010101000100","001100100010","010000110011","011001010101","001100110011","001100100010","001100100010","001100100010","010000110011","100110001001","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001100100001","001100100001","001000100010","001100110011","011001010101","011001010110","011001010101","010101000100","001100100010","010101000100","011101100111","001100110011","001100100010","001100100010","001100100010","010000110011","100001111000","100001111000","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001100100010","001100100010","001000100001","001000100010","001100100010","010101000100","011001010101","011001010110","010101000100","001000100010","010101000101","100001100111","001100110011","001100100010","001100100010","001100100010","001100110011","100001111000","100110001001","100001111001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100010","010101000100","010101010101","011001010101","010001000100","001000100010","010101000101","100001110111","001100110011","001100100010","001100100010","001000100010","001100100010","100001111000","100010001001","100001111000","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010000110011","010101000101","010101000101","010000110100","001000100010","010000110011","010101000101","001100100010","001100100010","001100100010","001000100010","001100100010","100001111000","100001111001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000101","010101000100","010000110011","001000100010","001100100011","010000110011","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000100","001100110011","001000100010","001100110011","010000110011","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010000110100","001100110011","001000100010","001100110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100010","010000110011","011001000100","011000110100","010000110011","010000110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","010101000100","100101111000","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000010001","001000010001","001100100010","010100110011","011101000100","011101000100","011101000100","011101000101","010000110011","010000110011","001000100010","001000100010","001000100010","001000100010","001000100001","010000110100","100101111001","100101111001","100110001001","100110001001","100010001001","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000010001","001000010001","001000100001","010100110011","011000110011","011101000100","011101000101","011101000101","011001000100","001100110011","010000110011","001000100010","001000100010","001000100010","001000100001","001000100001","010000110011","100101111000","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010100110011","011000110011","011101000100","011101000101","011101000101","010000110011","001100100010","010000110011","001000100010","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000101","011101100111","011101010110","100001100111","100001111000","100101111001"),
		("001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","011000110011","011000110011","011101000100","011101000101","011101000100","001100100010","001100100010","001100110011","001000100001","001000100001","001000100001","001000100001","001000100010","001000010001","000100010001","001000010001","010000100010","011000110011","011101000100","011101000101","011101010110"),
		("000100010001","001000010001","000100010001","000100010000","000100010000","001000010001","010100100010","011000110011","010100110011","010100110011","010000100010","001000100001","001100100010","001100100010","001000100001","001000100001","001000010001","001000100001","001000010001","000100010000","000100010000","001000010001","010000100010","011000110011","011000110011","011000110011","011101000100"),
		("000100010001","000100010001","001000010001","001000010001","001000010001","000100010000","001000010001","001000010001","001000100001","001000010001","000100010001","001000100001","001100100010","001100100010","001000100001","001000100001","001000010001","001000010001","000100010001","000100010000","000100010000","001000010001","010000100010","011000110011","011000110011","011000110011","011101000100"),
		("001000010001","001000010001","001000010001","001100100010","001000100010","001000010001","000100010000","000100010001","001000010001","001000100001","001000010001","001000100001","001100100011","001100100010","001100100010","010000110011","001100100010","001000100001","000100010000","000100010000","000100010000","000100010000","001000010001","010100100010","011000110011","011000110011","011101000101"),
		("001000010001","000100010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","000100010001","001000100001","001100110010","001100100010","001000010001","001000010001","011001010110","011101100111","010101000100","001100110010","001000100001","000100010001","000100010000","001000010001","001100100010","011001010101","100001111000"),
		("001000010001","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001100110010","001100100010","001000010001","001000010001","011001010101","100110001001","100110001001","100110001001","100001111000","011101100111","011001010110","010101010101","011001100110","100001111001","100010001001"),
		("001000010001","000100010001","000100010001","000100010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","001000100010","001000100001","001100110010","001100100010","001000010001","001000010001","010101000100","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001100100010","001000100001","001100110011","001100100010","001000010001","000100010001","001100110011","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100101111001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","001100110011","001000100001","001100110011","001100100010","001000010001","001000010001","001100100010","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","010000110011","001000100010","001100100011","001100100010","001000100001","001000100001","001000100010","100001110111","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000010001","000100010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010000","001000100001","010000110011","001100100010","001100110011","001100100010","001000100010","001000100010","001000100001","011101100111","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001","100110001001","100010001001","100010001001"),
		("001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000100010","010001000100","001100100010","001100100010","001100100010","001000100010","001000100010","001000100001","011001010110","100010001001","100001111001","100001111001","100001111001","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010101000100","010000110011","001100100010","001100100010","001000100001","001000100010","001000100001","010101000101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","000100010001","001000100010","010101000100","010000110011","001100100010","001000100010","001000100010","001000100001","001000100001","010000110011","011101100111","011101100111","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 27
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100010001001","100101111000","100101110111","100001100110","100001100110","100101110111","100001100111","100110001001","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110001011","100110001010","100101110111","100101010101","100001000100","011000110010","010100100001","010100100010","010100110010","011101000100","100101111000","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001010","100110011011","101010001001","100101100101","011000110011","010100100010","010000100010","010000100001","010000100001","010000100001","010100100010","011101000100","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010011010","100001010101","011000110010","010100100010","010000100001","010000100001","010000100001","010000100001","010000100001","010000100001","011101010101","101010011010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","100101111000","010100100010","010000100001","010000100001","010100100001","010100110010","011000110011","011001000100","011001000100","011101000100","100110001001","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100001010110","010100100001","010000100001","010000100001","010100100010","011101000100","100001010101","100101100110","100101100111","100101100111","100110001001","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110011010","100001111001","100001111001","100010001001"),
		("101110101100","101010101100","100110001010","011101010110","010000100001","010000100001","010000100001","011000110011","011101000101","100001010101","100101100110","100101100111","100101100111","100110001001","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","100110011010","011101010101","010000100001","010000100001","010000100010","011000110011","011101000101","100001000101","100001010101","100001010101","100001010110","100101100111","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101010101100","011101000101","010100100010","010100110010","010100100010","011000110100","011101000101","100001010101","100001010101","100001010110","100001010101","100001100111","100110001001","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","100101111000","011101000100","011101000100","011101000100","011101000100","011101000100","100001010101","100101010110","100101100110","100001010101","100101111000","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","101010011011","100001000101","011101000100","011101000100","011101000100","011101000100","011101000101","100001010110","100001010110","100001000101","100101111000","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101010101100","101010011100","101010011011","101110101100","100001100111","011101000100","011101000100","011101000100","011101000100","011101000100","100001010101","100001010110","100001010110","100110001001","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011011","101010011100","100110011011","101010101100","100110001001","011101000101","011101000100","011101000100","011101000100","011101000100","100001010101","100001010101","100001010110","100110001001","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("100110001010","101010011011","100110001010","100110001001","100101110111","011101000100","011101000100","011101000101","011101000101","011101000100","011101000101","100001010101","100001100111","100001111000","100110011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100010001001","100110001001","100101111000","011101000101","011101010101","011101000100","011101000100","011101000100","011101000101","011101000100","100001010101","100101111000","100101111001","100001111000","100110001001","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100001111000","011101100111","010100110011","001100100010","011101010101","011101000100","011101000100","011101000101","100001000101","100001010101","100001100111","100001111000","100001111000","100001111000","100001111000","100010001001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("010000110011","001100100010","001000100010","001000100001","011001010110","100001010110","011101000100","100001000101","100001010110","100001010101","100001100111","011001010110","011001000100","011001010101","011101100111","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100001","010101000100","100001111000","011101000101","100001010101","100001010110","011101000100","100001111000","011101100111","010101000101","011001010101","010101000100","010000110011","011101100110","100110001001","101010011010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("001000100010","001000100010","001100100010","001000100001","010101000100","100001111001","100001111000","100001010110","100001000101","011101000101","100110001010","011101100111","010101000101","011001010101","010000110100","001100100010","001100100010","010000110011","100001111000","101010011010","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001000100010","010000110011","100001111001","100010001001","100001111000","100001010110","100001111000","100110001010","011001010101","010101000100","011001010101","010000110011","001100100010","001100100010","001000100010","010101000100","101010011010","101010011010","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001000100010","001000100010","001000100010","001100100010","010101000100","011001010110","011001010110","011001010110","011101100111","011101100111","001100100010","010001000100","010101000101","001100100011","001100100010","001100100010","001100100010","010000110011","100110001001","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001100100001","001100100001","001000100010","010101000101","011001010110","011001010101","011001010101","010101000100","001100100010","010101000101","011001010110","001100100010","001100100010","001100100010","001100100010","001100100011","100001111000","100001111000","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001100100010","001100100010","001000100001","001000100010","010000110100","011001010101","011001010110","011001010101","010000110100","001000100010","011001010110","011101100110","001100100010","001100100010","001100100010","001100100010","001100100010","011101100111","100110001001","100001111001","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","010000110011","010101000101","011001010101","011001010101","010000110011","001000100010","011001010110","011101010110","001100100010","001100100010","001100100010","001100100010","001000100010","011101100111","100110001001","100001111000","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010101010101","011001010101","010000110011","001000100010","010000110100","010101000100","001100100010","001100100010","001100100010","001100100010","001000100010","011101100110","100001111001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010001000100","010101000100","010101010101","010000110011","001000100010","001100110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000100","001100110011","001000100010","010000110011","010000110011","001000100010","001000100010","001000100010","001100100010","001000100010","011001010110","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","010101000100","001100110011","001000100010","010000110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","010101010101","100110001001","100110001001","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110100","010000110011","001100100010","001000100010","010000110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100001","010001000100","100101111000","100110001001","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001100110011","010000110011","001100100010","001000100010","001100110011","001100110011","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100101111000","100101111001","100110001001","100110001001","100010001001","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000010001","001000010001","001000010001","001000100010","001100100010","010000110011","010101000100","010000110011","001000100010","001100110011","001100110011","001000100010","001000100010","001000100010","001000100001","001000100001","001100100010","100001111000","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","010000110011","011000110100","011101000100","011101000101","011101000100","010000110011","001100110011","001100110011","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","100001100111","100110001001","100110001001","100110001001","100110001001","100010001001","100101111001"),
		("001000010001","001000010001","001000010001","001000010001","000100010000","010000100010","011000110011","011101000100","011101000101","011101000101","011101000100","001100100010","001100110010","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","100001111000","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("000100010001","001000010001","000100010001","000100010000","000100010001","010100110011","011000110011","011101000100","011101000100","011101000100","010100110011","001000100001","001100110011","001100100010","001000100001","001000100001","001000010001","001000100001","001000010001","001000010001","010101000101","100001111000","100110001001","100101111001","100110001001","100110001001","100010001001"),
		("000100010001","000100010001","001000010001","001000010001","000100010001","010100100011","011000110011","011100110100","011101000100","011101000101","010000100010","001000100001","001100110011","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","000100010000","000100010000","001100100010","011001000100","011101000100","011101010110","100001010110","100001111000"),
		("001000010001","001000010001","000100010001","001000010001","001000010001","010000100010","011000110011","011000110011","011101000100","011000110011","001000100001","001000100001","001100110011","001100100010","001000010001","001000100001","001000010001","000100010001","000100010001","000100010000","000100010000","001000010001","010100100010","011000110011","011000110011","011000110011","011101000101"),
		("001000010001","000100010001","000100010001","001000010001","001000010001","001000100001","001100100001","001100100001","001100100010","001000100001","000100010001","001000010001","001100110011","001100100010","001000010001","001000010001","000100010001","000100010000","000100010001","000100010001","000100010001","001000100001","010100100010","011000110011","011000110011","011000110011","011101000100"),
		("001000010001","000100010000","001100100010","001100100010","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","000100010001","001000010001","001100110011","001100100010","001000010001","001000100001","001100100010","001000010001","000100010000","000100010000","000100010000","001000010001","010100100010","011000110011","011000110011","011000110011","011101000101"),
		("001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","001100100010","001100110011","001100100010","001000010001","001000010001","011001010101","011101100110","001100110010","000100010000","000100010000","000100010000","001100100001","010100100010","011000110011","011100110100","100001100110"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001100100011","001100110011","001100100010","001000010001","000100010001","010101000100","100110001001","100010001001","011001010110","001100110010","000100010001","000100010000","000100010001","011001000101","100001111000","100001111000"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","000100010000","001000100001","001100110011","010000110011","001100100010","001000010001","001000010001","001000100001","011101100111","100110001001","100110001001","100001111001","011101100111","010001000100","010000110011","100001111000","100110001001","100001111001"),
		("001000010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","010000110011","010000110011","001100100010","001000010001","001000010001","000100010000","011001010110","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000010001","000100010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010001","001000010001","001000010001","010000110011","010000110011","001000100010","001000010001","001000010001","001000010001","010101010101","100110001001","100110001001","100110001001","100110001001","100010001001","100010001001","100110001001","100010001001","100010001001"),
		("001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","000100010001","001000010001","010000110011","010000110011","001100100010","001000100010","001000100001","001000010001","010101000100","100010001001","100001111001","100001111001","100001111001","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000010001","010000110011","010000110011","001100100010","001000100001","001000100001","001000100001","010000110011","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010001","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010000","001000010001","010000110011","010000110011","001000100010","001000100001","001000100001","001000100001","001100100010","011101100110","011101100111","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 28
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100010001001","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","100010001001","100110001010","100010001001","100010001001","100010001001","100001111001","100110001001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001010","100110011011","101010011011","100110001001","100101111000","100110001001","100101111000","100101111000","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010011011","101010011010","100101100110","100001010100","100001000100","011100110011","011100110011","011101010101","100101111000","100110001010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011010","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010011011","100101110111","011000110010","010100100010","010100100010","010100100010","010100100010","010100100010","011101000100","100110001001","101010011010","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100101111000","100101010101","010100110010","010000100001","010000100001","010000100001","010000100001","010100100010","010100100010","100001100110","101010011011","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101100","101010101100","100110001010","100001010110","011000110011","010100100010","010100100010","010100110011","011000110011","011101000100","011101000101","011000110011","011101000101","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","100110011011","100001100111","010100100010","011101000100","100001010101","100001010110","100101100110","100101100111","100101100111","100001010110","011101000100","100110001010","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101110101100","100001100111","011000110010","100001000101","100001010101","100001010101","100101100110","100101100110","100101100110","100101100110","011101000101","100101111000","100110001001","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010101100","101010101100","100101111000","011000110011","011101000101","011101000100","011101000100","100001010101","100001010110","100001010101","100001010110","100001100110","100101111001","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110101101","101010101100","101010011100","101010001010","011101000100","011101000100","011101000100","011101000100","011101000101","100001010101","100001010101","100001010101","100101100111","100110001010","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101010101100","101010011100","101010011011","100101111000","011101000100","011101000100","011101000100","011101000100","011101000100","100001010110","100101100110","100001010110","100101100111","100110001010","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011011","101010011100","101010011011","100110001001","100001000100","011101000100","011101000100","011101000100","011101000100","100001010101","100101100110","100001010110","100101111000","100110001001","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("100110001010","101010011011","100110001010","100110001010","100001100111","011101000101","011101000100","011101000101","011101000101","100001010110","100101100110","100001100110","100001111000","100001111000","100110011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100010001001","100110001001","100110001010","101010011010","100110001001","100001010110","011101000100","011101000101","011101000100","100001010101","100001010110","100101111000","100110001001","100001111000","100110001001","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100001111000","100001111001","101010011010","101010011011","100110001010","100001010110","011101000100","011101000100","011101000101","100001010110","100001010110","100101111000","100001111000","011101100111","100001111000","100001111001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100001111000","100001111001","100110001010","101010011010","100110001001","100001010101","011101000100","011101000100","011101000100","100001010101","100001010110","100001100111","011001010101","011001000101","011101100111","100001111001","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100001111001","100001111000","100110001001","100001111000","011001000100","011101010101","011101000100","011101000011","011101000100","100001000101","100001010110","100001100111","011001010101","011001010101","011101100110","011101100111","100001111000","100110001010","101010011010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110001010","100001111000","011001010101","010000100010","001100100010","011101010110","011101000100","011101000100","011101000100","011101000101","100001010101","100001100111","011001010110","011001010101","010101010101","001100100010","010000110011","010101010101","100001111000","101010011010","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("011101100110","010000110011","001000100010","001000100010","001000100010","011001100110","100001010110","011101000100","011101000101","011101000101","011101000100","100001111000","011001010110","010101000101","010101000101","001100100010","001100100010","001100100010","001100100010","010101000101","100110001001","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001100100010","001000100010","001000100010","001000100010","001000100010","010101010101","100110001001","011101010110","100001000101","011101000100","011101010101","100110001010","011101100111","011001010101","010000110011","001100100010","001100100010","001100100010","001100100010","001000100010","010101010101","100001111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("001000100010","001100100010","001100100010","001100100001","001000100001","010101000101","100010001001","100010001001","100001100111","011101010101","100001111000","100110001010","011001010101","011101100111","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","010000110011","100001111001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("001000100001","001000100010","001100100010","001100100010","001000100001","010000110011","100001111000","100001111000","011101100111","011101100110","011101100111","011001010110","010000110100","100001100111","010000110011","001100100010","001100100010","001100100010","001100100010","001100100010","001100110011","100001111000","100001111000","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100010","001000100001","001000100001","001000100010","001100110011","011001010101","011001010110","011001010101","011001010101","010000110100","010000110011","100001110111","001100110011","001100100010","001100100010","001100100010","001000100010","001000100010","001100100011","100001111000","100010001001","100001111001","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010","010101000100","011001010110","011001010110","011001010101","010000110011","001100100010","010101000101","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","011001010101","011001010101","011001010101","010000110011","001100100010","010000110011","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","011001010101","011001010101","010101000101","001100110011","001100100010","010000110100","001100100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100010","011101100111","100110001001","100110001001","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010101000101","011001010101","010101000100","001100110011","001100100010","010000110100","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010000110100","010101000101","010000110100","001100100010","001100100010","010101000100","010100110011","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","011001010101","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100110011","010101000100","010000110011","001100100010","010100110100","011001000100","011101010101","100001010101","011101000101","001100100010","001000100010","001000100010","001000100001","010101010101","100110001001","100110001001","100010001001","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100010","001000100001","001100100010","010000110011","010000110011","001100100010","011000110011","011001000100","011101000101","100001010101","100001010110","001100110011","001000100001","001000100010","001000100010","011001010110","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","001000100001","010000110011","010000110011","001100100010","010000110011","010101000100","011101000101","100001010101","100001010101","001100100010","001000100001","001000100001","001000100010","011101100111","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","001000100001","001000010001","001000010001","001100110010","010000110011","001000100010","001000100001","010000110100","011000110100","100001000101","011101000101","001100100010","001000100001","001000100010","001000100001","001100110011","100001111000","100110001001","100110001001","100110001001","100001111001"),
		("000100010001","001000010001","000100010001","000100010001","000100010001","001000100001","001000100001","001000010001","000100010001","001100100010","010000110011","001000100010","001000100001","001100110011","001000010001","010100110011","010100110011","001000100010","001000100010","001000100001","001000100001","001000010001","011101100110","100110001001","100110001001","100110001001","100001111001"),
		("000100010001","000100010001","001000010001","001000010001","000100010001","001000010001","001000100001","001000010001","000100010001","001000100001","010000110011","001000100010","001000100001","001100110010","000100010001","001000100001","001000100001","001000100001","001000100010","001000100010","001000100001","010101000101","100101111001","100010001001","100001111001","100001111001","100101111000"),
		("001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000100001","001100110011","001000100010","001000100010","001100100010","001000010001","001000100001","001000010001","001100100010","001000100010","001000100001","001100110011","100001111000","100110001001","100110001001","100001111001","100001111000","100001111000"),
		("001000010001","000100010001","000100010001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000100001","001100110011","001100100010","001100100010","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000100010","011001010110","100110001001","100110001001","100110001001","100010001001","100010001001","100001111000"),
		("000100010001","000100010000","000100010000","000100010000","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","001100100010","001100100010","001100110010","001000010001","001000010001","001000010001","001000100010","011001010101","100001111000","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("001100100010","001100100010","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001100100010","001000100010","001100100010","001100110011","001000010001","001000010001","010001000100","100001110111","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001"),
		("011101000101","011101000101","001100100010","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","001000100001","001000010001","010000110011","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("011101000100","011101000101","010100110011","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","000100010001","001000100001","001000100010","010000110011","001100110011","001000100010","001000100010","001100100010","011101100111","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100110001001","100001111001"),
		("011101000101","100001000101","011000110100","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","000100010001","001100110011","010101000100","010000110011","001100100010","001000100010","001000100010","001000100001","010101000100","100110001001","100110001001","100110001001","100110001001","100110001001","100010001001","100110001001","100110001001","100001111001"),
		("011101000100","100001000101","011001000100","001000100001","001000010001","001000010001","001000010001","000100010001","000100010001","000100010000","001100110010","010101000101","010101000100","010000110011","001000100010","001000100010","001000010001","001100110011","100001111001","100110001001","100110001001","100110001001","100010001001","100010001001","100110001001","100010001001","100010001001"),
		("011000110011","011101000100","011000110011","001000010001","000100010001","001000010001","001000010001","000100010001","001000010001","000100010000","001100100010","010101010101","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","011101100111","100010001001","100001111001","100001111001","100001111000","100001111001","100001111001","100001111001","100001111001"),
		("001000100001","001100100001","001100100001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000100010","010101010101","010101000100","010000110011","001100100010","001000100010","001000100010","001000100001","010101010101","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("000100010000","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010000","001000100001","010101000100","010101000100","010000110011","001100100010","001000100001","001000100001","001000100001","010000110011","011101100111","011101100111","011101100111","011101100110","011101100111","011101100111","011101100111","011101100111"))
	-- 29
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100010001001","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","100010001001","100110001010","100010001001","100001111001","100001111001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001010","100110011011","101010011011","100110001010","100110001010","100110001010","100010001001","100110001001","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010011011","101010101100","100110001010","100110001010","100110001010","101010011010","101010011011","101010011011","101010101100","101010011011","101010011010","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100110001010","101010011011","100101111000","100101100110","100001010101","100001010100","100001010101","100001100111","101010001001","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101100","101010101100","100110001010","101010011011","100101111000","100001000100","011101000011","011000110010","010100100010","010100100010","011000110011","011101000011","100001100110","101010011011","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","101010011011","101010101100","100101110111","011000110010","010000100010","010100100010","010100100010","010000100001","010100100010","010100100010","011000110011","100101111000","100110001010","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101010101100","101010101100","100101110111","011000110010","010100100010","010100100010","010100110011","011000110011","011101000100","011000110011","010100100010","100001010110","100110001010","101010011011","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010011100","101010101100","101010101100","100101100111","100001000100","100001000101","100001010101","100101010110","100101100110","100101100110","100001010101","010100100010","011101010110","101010011011","101010011100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110101101","101010101100","101010011011","101010101100","100001010101","100001010101","100001010101","100001010101","100001010110","100101010110","100101100110","100001010110","011000110011","011101010110","101010011011","101010011011","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101010101100","101010011100","101010011011","101010101100","100101100111","100001010101","011101000100","011101000101","100001010101","100001010101","100001010110","100001010110","011000110011","100001100111","101010011011","101010011011","101010011011","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010101100","101010011011","101010101100","101010001001","100001010101","011000110011","011101000100","100001010101","011101000100","011101000101","100001010110","011101000100","100001111000","101010011011","101010011011","101010011011","101010011011","101010011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("100110011011","101010011011","100110001010","101010011010","100101111001","100001010101","011101000100","011101000101","100101010110","100101100110","100101100110","100101010110","100001010110","100001100111","100110011010","101010011011","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100010001001","100110001001","101010011010","101010011010","100101100111","100001010101","011101000100","011101000100","100001010101","100101100110","100101100110","100101100110","100101100110","100001111000","100110001001","101010011010","101010011010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100110001001","101010011010","101010011011","100110001001","100001010110","011101000100","011101000100","100001010101","100101100110","100001100110","100001010110","100001100110","100001111000","100001111000","100001111001","100001111001","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100001111000","100001111001","100110001010","101010011010","100110001010","100101100111","011101000100","011101000011","011101000100","100001010110","100001010110","100001010110","011001010101","011001010101","100001111000","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110001010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100001111001","100001111000","100110001001","101010011011","100110001010","100101111000","100001000101","011100110011","100001000101","100001010110","100001010110","011101010101","011001010101","011001010101","100110001001","100001111001","100001111001","100110001010","100110001010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110001010","100001111000","100110001001","101010011011","100110001010","100101111000","100001010101","011101000100","011101000100","100001000101","100001010110","011101010101","010101000101","011001010101","100110001001","100001111001","100001111001","100110001010","100110001010","101010011010","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("101010011010","100110001001","100001111001","101010011010","100110001001","100001111000","100001010101","011101000100","011100110100","011101000100","100001010101","011101010101","010101000100","011001010101","011001010110","011101100111","100001111000","100001111001","100110001010","101010011010","101010011010","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100001111001","100110001001","011101100110","011001000100","100001010101","011101000100","011100110011","011101000100","100001010110","100001010101","011001010101","010101000101","001100100010","001100100010","001100110011","010000110100","011001010101","011101100111","100001111001","100001111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("100110001001","100101111000","011101100111","010100110011","001100100001","010000110011","100001100111","011101000100","011101000100","011101000100","100001000101","011101000101","011101100111","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","010000110011","010101010101","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100001100111","011001000100","001100100010","001000100001","001000100001","001100100010","100001111000","100001100110","011101000100","011101000101","011101000100","011101010110","100001111001","011001010101","001100100010","001100100010","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","011001010101","100001111001","100010001001","100001111001","100001111000"),
		("010000110011","001000100010","001000100010","001000100001","001000100001","001100100010","011101100111","100010001001","100001100111","011101000101","011101000101","100001111000","100110001001","011001010101","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","010000110011","100001111000","100010001001","100001111001","100001111000"),
		("001000100001","001000100010","001000100001","001000100001","001000100001","001000100010","011101100110","100001111001","100001111000","011101010110","011101100111","100010001001","100001111000","010001000100","001100100010","001100100010","001100100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100001111001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000100","010101000100","010101000101","011001010110","011001010101","001100100011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100110001001","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101010101","011001010101","011001010101","011001010101","010101000101","001100110011","001000100010","001000100010","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","010101000101","100110001001","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001100100010","010101000100","011001010101","011001010101","010101010101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010000110100","100110001001","100001111001","100001111000"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","010001000100","011001010101","011001010101","010101000101","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001100110011","100001111000","100001111001","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","011001010101","010101010101","010101000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100010001001","100001111000"),
		("001000010001","001000010001","001000100001","001000100001","001000100010","001000100001","001000100010","001000100001","001100100010","010101000101","010101000101","010001000100","010101000100","001100100011","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","011101100111","100110001001","100001111001"),
		("001000100001","001000010001","001000010001","001000100001","001000100010","001000100001","001000100001","001000010001","001000100001","010101000100","010101000100","010001000100","010101000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100001","011001010110","100110001001","100001111001"),
		("010100100010","001000010001","001000010001","001000010001","001000100010","001000100010","001000100001","001000010001","001000100001","010000110100","010101000100","010000110100","010001000100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100001","011001010101","100110001001","100001111001"),
		("011101000100","010000100010","000100010001","000100010001","001000100001","001000100001","001000100001","001000010001","001000010001","001100110011","010101000100","010001000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001100100010","001000100010","001000100001","001100110011","011101100111","100010001001"),
		("100001010101","011000110100","001000100001","000100010001","001000010001","001000100001","001000100001","001000010001","001000010001","001100100010","010000110100","010000110100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","011000110011","010100110011","010000100010","001000100001","001100110011","100001111000"),
		("100001010110","100001000101","001100100010","000100010001","001000010001","001000100001","001000010001","001000010001","001000100001","001000100010","010000110011","010000110100","010000110100","001100100010","001000100001","001000100001","001000100001","001000100001","001000100010","001000100010","001100100010","011000110100","011101000101","100001010101","010100110011","010101000100","100001111000"),
		("100001010101","100001010101","010000100010","000100010000","001000010001","001000010001","001000100001","001000010001","001000100001","001000100001","010000110011","010000110100","010000110100","001100110011","001000100001","001000100001","001000100010","001000100010","001000100001","001100100010","010100110011","011101000100","011101000101","100001010101","011101000101","011101100111","100001111001"),
		("100001010101","100001010110","010000100010","000100010000","001000010001","001000010001","001000010001","001000100001","001000010001","001000010001","001100110011","010000110011","010000110011","010000110011","001000100001","001000010001","001000100001","001000100001","001000100001","001100100001","010100110011","011101000100","011101000101","100001010101","100001010101","100001111000","100010001001"),
		("100001000101","011101000101","001100100001","000100010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","010000110011","010000110011","001000100001","001000010001","001000010001","001000010001","000100010000","000100010000","001100100001","010100110011","011101000100","100001010101","011101000101","100001100111","100110001001"),
		("010000100010","001100100001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010101000100","010000110100","010000110100","001100100010","001000100001","001000010001","000100010000","000100010000","000100010000","000100010000","001000100001","010100110011","011000110100","011001000100","100001111000","100010001001"),
		("001000010001","000100010001","000100010000","001000010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000010001","001000100001","010000110011","010000110100","010000110011","001100100010","001000100001","000100010001","001000010001","001000100001","000100010000","001000100001","001000010001","001000010001","001100100001","011001010110","100110001001","100001111001"),
		("001100100010","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","001000100001","001100100010","010000110011","001100110011","001100100010","001000100001","001000010001","001000010001","001000100001","000100010000","010101000100","011001010110","001100110011","010101000101","100001111000","100110001001","100001111001"),
		("100001110111","011001010101","001000100001","000100010001","001000010001","001000010001","001000010001","000100010001","000100010001","001000010001","000100010001","001100100010","010000110011","010000110011","001100110011","001000100010","001000100001","001000100001","001000100001","001000010001","010001000100","100110001001","100001111000","100001111000","100110001001","100010001001","100010001001"),
		("011101100111","001100110011","001000010001","000100010001","000100010001","001000010001","001000010001","000100010001","001000010001","000100010001","001000010001","010000110011","010101000100","010101000100","010101000100","010000110100","001000100010","001000100001","001000100001","001000100001","001100110011","100001111000","100001111001","100001111001","100001111001","100001111001","100001111001"),
		("011001010110","001100100010","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","001000010001","000100010000","001000010001","010101000101","010101000101","011001010101","011001010110","010101000100","001100100010","001000010001","001000010001","001000100001","001000100010","011001010110","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("010000110011","001000010001","001000010001","001000010001","001000010001","001000010001","000100010001","001000010001","001000010001","000100010000","000100010001","010001000100","010101000100","010101000101","010101010101","010101000100","010000110011","001000100001","001000010001","001000010001","001000100001","010101000101","011101100111","011101100111","011101100111","011101100111","011101100111"))
	-- 30
	,

		(	("100110011011","101010011011","101010011011","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111001","100001111000","100001111000","100110001010","100110011010","100110011010","100110001010","100001111001","100010001001","100010001001","100001111000","100001111000","100001111000","100001111000","100001111000","100001111000"),
		("101010101100","101010101100","101010101100","101110101100","101010011011","100010001010","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100010001001","100110001010","100110001010","100010001001","100001111000","100001111000","100001111001"),
		("101110101100","101110101100","101110101100","101010101100","100110011011","100010001001","100001111001","100001111001","100110001010","100110001010","100110001010","100001111001","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110011010","100110001010","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101110101101","101010011011","100110001010","100110001010","100110001010","100010001001","100110001010","100010001001","100001111001","100001111001","100001111001","100110001001","100110011010","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","100110001010","100001111001","100001111001","100001111001","100001111001"),
		("101010011100","101010011011","100110001010","100110011011","101010011011","100110001010","100110001010","100110001010","100010001001","100110001001","100110001010","100110001010","100010001001","100110001001","101010011011","101010101100","101010101100","101010011011","100110001001","100110001001","100110001010","100110001001","100001111001","100010001010","100110001010","100001111001","100010001001"),
		("100110011011","100110001011","100110011011","101010011011","101010011011","100110001010","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","100110001010","100110001001","100110001010","101010101100","101010101100","101010011011","100110001010","101010011011","101010011011","101010011011","100110001010","100001111001","100010001001","100001111001","100010001001"),
		("101110101100","101010101100","100110011011","101010011011","101010101100","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","101010101100","101010011011","101010011010","100110001010","100110001010","100110001010","100110001010","101010011011","101010101100","101010011011","101010011011","101010011011","100110001001","100001111001","100001111001","100010001001"),
		("101110101100","101110101101","101010011011","100110001010","101010011011","100110001010","100110001010","100110001010","101010011011","101010011011","101010011011","101010101100","101010011011","101010011011","101010011011","100110001010","100110001001","101010011011","101010011100","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100010001001"),
		("101110101100","101010101100","100110001010","101010011011","100110001010","100110001010","100110001010","100110011010","101010001001","100101110111","100101100111","100101100110","100101110111","101010001010","101010011011","100110001010","100110001010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","101010011011","101010101100","101010011011","100110001010","100110001010","100101110111","100001010100","100001000011","011000110010","010100100010","010100100010","011101000100","100101100111","100110001001","100110001001","101010011010","101010011011","101010011011","101010011011","101010011011","101010011011","101010011011","100010001001","100001111001","100001111001"),
		("101010011011","100110011011","101110101100","101110101101","101010101100","100110001010","100110001010","100001010101","010100100010","010100100010","010100100010","010100100010","010100100010","010100100010","011000110011","100001100111","101010011010","100010001001","100010001001","100110011010","101010011011","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101110101101","101010011100","101010101100","101110101101","101010101100","100110001010","100101111000","100001000100","010100100010","010000100001","010100100010","010100110010","011000110011","011000110011","010100100010","011101000100","101010011011","100110001010","100001111001","100001111001","100110011010","101010011011","100110001010","100001111001","100010001001","100001111001","100001111001"),
		("101110111101","101010101100","101010011011","101110101100","101010101100","100110001010","100101111000","100001010100","011101000100","011101000101","100001010101","100001010110","100101100110","100101100110","011000110011","011001000100","101010011011","101010011010","100110001010","100001111001","100001111001","100010001001","100001111001","100010001001","100110001010","100001111001","100001111001"),
		("101110101100","101010101100","101010011011","101110101100","101010011100","100110001010","100001100111","100001000100","100001010101","100001010110","100001010110","100001010110","100101100110","100101100110","011101000101","011000110011","100110001010","101010011010","101010011010","100110001010","100001111001","100110001010","100010001010","100001111001","100001111001","100001111001","100001111001"),
		("101010101100","101010101100","101010011011","101010101100","101010011011","100110001010","100001100111","011101000100","100001000101","011101000101","100001010101","100001010101","100001010110","100101100110","100001010101","011001000100","101010011010","101010011011","101010011010","100110001010","100010001001","101010011011","101010011011","100110001010","100001111001","100001111001","100001111001"),
		("101010011011","101010011011","100110001010","101010011010","101010011011","100110001010","100101111000","100001010101","011101000100","011000110011","011101000101","100001010101","011101000100","100001010101","100001010101","011101010110","101010011011","101010011010","100001111001","100001111000","100001111001","100110001010","101010011011","101010011010","100110001001","100001111001","100001111001"),
		("100010001001","100110001010","101010011010","101010011010","100110001010","100110001010","100101111001","100101100111","011101000100","011101000100","011101000101","100101100110","100001010110","100101100110","100101010110","100001010110","100110001010","100110001001","100001111000","100110001010","100110011010","100001111001","100110001010","101010011011","100110001010","100001111001","100001111000"),
		("100001111001","100110001001","101010011010","101010011011","100110011010","100110001010","100101111000","100101100110","100001000101","011101000100","011101000101","100001010110","100001100110","100001100111","100001100110","100001100110","100001111000","100001111000","100110001001","101010011011","101010011011","100110001001","100010001001","101010011010","100010001001","100001111000","100001111000"),
		("100001111000","100010001001","101010011010","101010011010","100110001010","100110001001","100101111001","100101100111","100001010101","011101000100","011101000100","100001010110","011101010101","011001010101","011101010110","100001111000","100001111001","100110001010","101010011010","101010011011","101010011011","100110011010","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100001111001","100001111000","100110001010","101010011011","100110001010","100101111001","100110001001","100110001001","100001010110","011101000100","011100110100","011101000101","011001010101","011001010101","100001111000","100001111001","100010001001","100110001010","100110001010","101010011011","101010011011","101010011011","100110001001","100001111000","100001111000","100001111000","100001111000"),
		("100110001010","100001111000","100110001001","101010011011","100110001010","100001111000","100110001001","100110001010","100001100111","011101000100","011101000100","100001010101","011001010101","011001010101","100001111000","100001111001","100001111001","100110001010","100110001010","101010011010","101010011011","101010011011","100110001001","100110001001","100110001001","100001111000","100001111000"),
		("101010011010","100110001001","100001111001","101010011010","100110001001","100001111001","100001111001","100110001001","100001100111","011101000100","011101000100","011101000101","011001000101","010101000101","100001110111","100001111001","100001111000","100001111001","100110001001","100110001010","101010011010","100101111001","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("101010011011","100110001001","100001111001","100110001010","100110001010","100001111001","100001111000","100110001001","100001010110","011100110011","011100110011","011101000100","011101010101","011001010110","100001100111","011101100111","100001111001","100001111001","100001111001","100110001010","100110001001","100001111000","100001111000","100110001001","100110001001","100001111000","100001111000"),
		("100110001001","100101111001","100110001001","100110001001","100110001001","100001111000","100001100111","100001100111","100001010101","011101000100","011100110100","011101000101","100001100111","011101100111","100001100111","010101000100","010101000100","011101100111","100001111000","100010001001","100001111001","100110001001","100001111000","100001111001","100001111001","100001111000","100001111000"),
		("100101111000","100101111000","100110001001","100001111000","100001100110","011001000100","010100110011","011101010101","100001010110","011101000100","011101000100","011101000100","100001100111","011101100111","100001100111","010101000101","001000100010","001100100010","010000110100","011001010110","100001111000","100110001001","100001111001","100001111000","100010001001","100001111001","100001111000"),
		("100110001001","100110001001","100001100110","011001000100","001100100010","001000100001","001000100001","011001000101","100101111000","011101000100","011101000100","011101000100","100001100111","100001111000","100001111001","010101000101","001000100010","001100100010","001000100010","001000100010","001100100010","010001000100","011101100111","100001111000","100010001001","100001111001","100001111000"),
		("100001100110","011001000100","001100100010","001000100001","001000100001","001000100001","001000100001","011001010101","100110001001","100001100111","011101000101","011101000100","011101010101","100001100111","100110001001","010001000100","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001100100010","010000110100","011101100111","100001111001","100001111000"),
		("001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","011001010101","100001111000","100010001001","100001100110","011101010101","011101100111","011101100111","100001110111","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","010101000100","100001111001","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","010000110011","010101000100","010101000101","011001010101","011101100111","011101100111","011101100110","010101000101","001000100010","001000100010","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100110011","100001111000","100001111000"),
		("001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000100","010101000100","011001010101","010101000101","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100010","100001111000","100001111001"),
		("001000100001","001000010001","001000100001","001000100001","001000010001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000101","010101000101","010101000101","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111","100001111001"),
		("001000100001","001000010001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100010","010101000100","010101000101","010101000101","010101000101","010101000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010101010101","100110001001"),
		("001000010001","001000010001","001000100001","001000100001","001000100001","001000100001","010000110011","011001000100","010101000100","010101000100","010101000101","010101000101","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","010000110100","100110001001"),
		("001000010001","001000010001","001000010001","001000100001","001100100010","011001000100","011101000101","011101000100","011000110011","010100110100","010101010101","010101000100","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001100100011","100001111000"),
		("001000100001","001000010001","000100010001","001000010001","011001000100","011101000100","011000110100","011000110100","010100110010","010000110011","011001010101","010101000100","010101000100","010101000100","010000110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011101100111"),
		("001000100001","001000010001","000100010001","001000100001","011101000100","011101000100","011101000100","011101000100","011101000101","011001000100","010101000101","010101000100","010101000100","010101000100","010000110011","001100100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","011001010110"),
		("001000100001","001000010001","001000010001","001100100001","011000110100","011101000101","011101000101","011101000101","010100110011","001100100010","010001000100","010101000100","010001000100","010001000100","001100110011","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100010","001000100010","001000100010","010001000100"),
		("001000100001","001000100001","001000100010","001100100010","011000110100","011101000101","011101000100","011001000100","001100100010","001000100001","001100110011","010000110100","010001000100","010000110100","001100100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100010","001000100001","001000100001","001000100010","001000100010","001100100010"),
		("001100100010","001100100010","001000100001","001100100010","011000110011","010100110011","001100100001","001000010001","001000100001","001000100001","001100100011","010000110011","010001000100","010001000100","010000110011","001100100010","001000100010","001000100001","001000100001","001000100001","001000100010","001000100010","001000100001","001000100001","001000100001","001000100001","001000100010"),
		("001000100010","001000100010","001000100001","001100100001","010000100010","001100100001","000100010001","001000100001","001000100001","001000100001","001100100010","010000110011","010001000100","010000110100","010000110011","001100100010","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000100001","001000100001"),
		("001000100001","001000100010","001100100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","010000110100","010000110100","010000110011","001100100010","001000100001","001000100001","001000100010","001000100001","001000100001","001000100001","001000100001","001000010001","001000010001","001000010001","001000100001"),
		("001000100001","001000100010","001100100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001","001100100010","010000110011","010000110011","010000110100","010000110011","001100110011","001000100001","001000010001","001000100010","001000100010","001000100010","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001"),
		("001000100001","001000010001","001000010001","000100010001","001000010001","001000010001","001000010001","000100010001","001000100001","001000100001","001100100010","010000110011","010000110011","010000110100","010000110011","001100110011","001000100010","001000010001","001000100001","001000100010","001000100001","001000100001","001000010001","001000010001","001000010001","001000010001","001000010001"),
		("001000100001","001000100001","001000100001","001100100010","001000010001","001000010001","001000010001","000100010001","001000010001","001000100001","001000100010","010000110011","010000110011","010000110011","010000110011","010000110011","001000100010","001000010001","001000010001","001000100001","001000100001","001000100001","001000010001","000100010001","000100010001","001000010001","001000010001"),
		("011101100110","011001010110","011101100111","011101010110","001000010001","001000010001","001000010001","000100010000","001000010001","001000100001","001000100010","010000110011","010000110011","010000110011","010000110011","001100110011","001100100010","001000100001","001000100001","001000100001","001000100001","001000010001","000100010001","000100010000","000100010000","000100010001","001000100001"),
		("100001111000","100001111000","100001111000","010101000101","001000010001","001000010001","001000010001","000100010001","001000010001","001000100010","001000100010","001100100010","010000110011","010000110011","001100110011","010000110011","001100110011","001100100010","001000100010","001000100001","001000100001","000100010001","000100010000","000100010000","000100010000","001000010001","010000100010"),
		("100001110111","100001111000","100001111000","010000110011","000100010001","001000010001","001000010001","001000010001","001000010001","001000100001","001000100001","001000010001","001100100010","010000110011","010000110011","010101000100","010101000100","010000110011","001000100010","001000010001","001000010001","000100010001","000100010000","000100010000","000100010000","001000010001","010000100010"),
		("011101100111","011101100111","011101100110","001100100010","000100010001","001000010001","000100010001","001000010001","001000010001","001000010001","001000100001","001100100010","010000110011","010101000100","010101010101","010101010101","010101010101","010000110100","001100100010","001000010001","001000010001","000100010001","000100010000","000100010001","001000100001","001000010001","010000100010"))
	-- 31

	);

    type color_sprite is array (0 to 15, 0 to 15) of std_logic_vector(0 to 11);

    constant BRICK_ROM : color_sprite := (
        ("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
        ("000000000000","000100000000","001100000000","001100000000","001100000000","001100000000","001100000000","000000000000","001100000000","001100000000","001100000000","001100000000","001100000000","001100000000","001000000000","000000000000"),
        ("000000000000","001100000000","110000010000","101100010000","101100010000","101100010000","101000010000","001000000000","101000010000","101100010000","101100010000","101100010000","101100010000","101100010000","001100000000","000000000000"),
        ("000000000000","010000000000","110100010000","110100010000","110100010000","110100010000","101000010000","001000000000","101100010000","110100010000","110100010000","110100010000","110100010000","101100010000","001100000000","000000000000"),
        ("000000000000","010000000000","110100010000","110100010000","110100010000","110100010000","101000010000","001000000000","101100010000","110100010000","110100010000","110100010000","110100010000","101100010000","001100000000","000000000000"),
        ("000000000000","000100000000","001100000000","001100000000","001100000000","001100000000","001000000000","000000000000","001100000000","001100000000","001100000000","001100000000","001100000000","001100000000","000000000000","000000000000"),
        ("000000000000","001100000000","101100010000","100100010000","001000000000","011000000000","101100010000","101000010000","101000010000","101000010000","010100000000","001100000000","101100010000","100100010000","001000000000","000000000000"),
        ("000000000000","010000000000","111000010000","110000010000","001100000000","100000010000","111000010000","111000010000","111000010000","110100010000","011100000000","010000000000","111000010000","110000010000","001100000000","000000000000"),
        ("000000000000","001100000000","101100010000","100100010000","001000000000","011000000000","101100010000","101100010000","101100010000","101000010000","010100000000","001100000000","101100010000","100100010000","001000000000","000000000000"),
        ("000000000000","000100000000","001100000000","001100000000","001100000000","001100000000","001100000000","001000000000","000000000000","001100000000","001100000000","001100000000","001100000000","001000000000","000000000000","000000000000"),
        ("000000000000","010000000000","111000010000","110100010000","110100010000","110100010000","110100010000","100100010000","001000000000","110000010000","111000010000","110100010000","111000010000","110000010000","001100000000","000000000000"),
        ("000000000000","001000000000","011100010000","011100010000","100000010000","011100010000","011100010000","010100000000","000000000000","011100000000","100000010000","100000010000","011100010000","011000000000","001000000000","000000000000"),
        ("000000000000","000100000000","011000000000","010100000000","000100000000","001100000000","011000000000","011000000000","011000000000","010100000000","001000000000","000100000000","011000000000","010100000000","000100000000","000000000000"),
        ("000000000000","010000000000","111000010000","110000010000","001100000000","100100010000","111000010000","111000010000","111000010000","111000010000","011100000000","010000000000","111000010000","110000010000","001100000000","000000000000"),
        ("000000000000","001000000000","010000000000","010000000000","000100000000","001000000000","010000000000","010000000000","010000000000","010000000000","001000000000","000100000000","010000000000","010000000000","001000000000","000000000000"),
        ("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000")
    );
    
	type apple_gif_sprite is array (0 to 1, 0 to 15, 0 to 15) of std_logic_vector(0 to 11);
	constant apple_GIF_ROM : apple_gif_sprite := (

		(	("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","000000000000","110010100010","000000000000","000000000000"),
		("000000000000","111111000011","111111000011","110010100010","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111111000011","111111000011","110010100010","000000000000"),
		("000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","100001010011","000000000000","000000000000","110010100010","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","100001010011","011001110011","000000000000","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","000000000000","111001110110","111001100110","000000000000","100001010011","011101000010","011001100011","011001110011","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","111001110111","111001100110","110100110011","110100110011","011101000010","010001100010","010001100010","110000110010","110000110011","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","111001110111","111001100110","111000110011","111110101010","111000110011","110000100010","110000100010","110000100010","111000110011","110100100010","110000110011","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","111001100110","111001000100","111110101010","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","110100100010","101100110011","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","111001010101","111000110011","111110101010","111000110011","111000110011","111000110011","111000110011","111000110011","110100100010","110000110011","101000110011","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","110100110011","111000110011","111110011001","111000110011","111000110011","111000110011","110100100010","110000110011","101000110011","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","110000110011","110100100010","111000110011","111000110011","111000110011","110100100010","110000110011","101000100010","100000100010","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","110010100010","000000000000","110000110011","101100110011","100100100010","000000000000","110000110011","101000110011","100000100010","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","111111000011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","110010100010","000000000000"),
		("000000000000","000000000000","000000000000","110010100010","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000"))
	-- 0
	,

		(	("000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111010110011","011101110000","000000000000"),
		("000000000000","000000000000","000000000000","111010110011","111101110000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111111110111","111111010100","111010110011","101110010010","000000000000"),
		("000000000000","111111110000","111111000011","111010110011","101110010010","000000000000","000000000000","000000000000","000000000000","000000000000","100101000011","111011001000","111111010101","111111000011","111111000011","000000000000"),
		("000000000000","111111010011","111010110011","110110100010","011101110000","000000000000","000000000000","000000000000","000000000000","100001010011","100001010011","100101100100","111111010101","111111010011","111101110000","000000000000"),
		("000000000000","111111110000","111010110011","000000000000","000000000000","111001100110","111001100110","000011111111","100001000011","100001010011","011001110011","010101110011","000000000000","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","000000000000","111001110111","111001100110","111001100110","110001000100","100001010011","011101000011","011001100011","011001100011","100101010011","111111110000","111010110011","111101110000"),
		("000000000000","111010110011","101101110011","111001110111","111001110111","111001100110","111001010101","110100110011","100001000011","010101100010","011001100010","110000110011","110000110011","110101100011","111010110011","101110010010"),
		("111111010100","111010110011","110110000100","111001110111","111001100110","111001100110","111010001000","111000110011","110100110011","110100110011","110100110011","111000110011","111000110011","110000110011","110101110010","000000000000"),
		("111111010101","111010110010","111001100110","111001100110","111001010101","111010011001","111001000100","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","101100110011","101100110011","111010110011"),
		("111111010100","111010110011","110101110100","111001010101","111001000100","111010011001","111001000100","111000110011","111000110011","111000110011","111000110011","110100110011","110000110011","101000100011","110110000011","111010110011"),
		("000000000000","111010110011","101101110011","110101010101","111000110011","111001000100","111001110111","111000110011","111000110011","111000110011","110100110011","110000110011","101000110011","101000100010","101101110011","111010110011"),
		("000000000000","000000000000","000000000000","101000100010","110000110011","111000110011","111000110011","110100110011","111000110011","110100110011","110000110011","101000100010","100100100010","011100100010","000000000000","000000000000"),
		("000000000000","000000000000","000000000000","111100000000","110101010011","110000110011","110000100010","101000100010","110000110011","110000110011","101000110011","100000100010","100000100011","000000000000","000000000000","000000000000"),
		("000000000000","000000000000","111111110000","111111000011","111010110011","110001100010","101100110011","100100100010","000000000000","110000100010","101000110011","100000100010","111111111111","111111010101","111111110011","111010110011"),
		("000000000000","000000000000","111111010011","111010110011","110110100010","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111111011001","111111010101","111111000010","111010110011"),
		("000000000000","000000000000","111111110111","111010110011","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","000000000000","111111110111","111111010110","111111000011","111010110010"))
	-- 1

	);

	type color_sprite_8 is array (0 to 7, 0 to 7) of std_logic_vector(0 to 11);
	constant SNAKE_ROM : color_sprite_8 := (
		("010101100010","011010000010","011010000010","011010000010","011010000010","011010000010","011010000010","001001010001"),
		("011010000010","010011000001","001110110001","001110110001","001110110001","001110110001","001110110001","001001100001"),
		("011010000010","001110110001","000110100001","000110100000","000110100000","000110100001","000110100000","001001100001"),
		("011010000010","001110110001","000101110001","001010100001","001010100001","001001110001","001010100001","001001100001"),
		("011010000010","001110110001","000110100001","001010010001","001010010001","001010100001","001010110000","001001100001"),
		("011010000010","001110110001","000110100001","001010100001","001010100001","001010100001","001010110000","001001100001"),
		("011010000010","001110110001","000110110000","001010110000","001010110000","001010110000","001010110000","001001100001"),
		("001001010001","001001100001","001001100001","001001100001","001001100001","001001100001","001001100001","000101010001")
	);

--    vgaRed <= COLOR_ROM(row, col)(11 downto 8);

    constant img_size_x : natural := 16;
    constant img_size_y : natural := 16;

    signal is_img_painted : std_logic;
    signal img_clr : std_logic_vector(11 downto 0);

    signal img_x : unsigned(10 downto 0) := to_unsigned(50, 11);
    signal img_y : unsigned(10 downto 0) := to_unsigned(50, 11);
    
    signal rgb : std_logic_vector(11 downto 0);
    
    signal current_frame_gif : unsigned(11 downto 0) := to_unsigned(0, 12);

    signal brick_clr : std_logic_vector(11 downto 0);

	signal snake_clr : std_logic_vector(11 downto 0); -- snake colour signal
begin
    led <= switch;
    start <= switch(7);
    
    process(pixel_clk)
    begin
        if rising_edge(pixel_clk)then
             if yCount = to_unsigned(1, yCount'length) and xCount = to_unsigned(1, xCount'length) then
                current_frame_gif <= current_frame_gif + 1;
             end if; 
        end if;
    end process;
    
    is_img_painted <= '1' when (xCount >= img_x and xCount < img_x + 16 and yCount >= img_y and yCount < img_y + 16) else '0';
    --is_img_painted <= '1';
--    img_clr <= ROM((yCount - img_y) mod img_size_y)((xCount - img_x) mod img_size_x) when is_img_painted = '1' else '0';
--    img_clr <= COLOR_ROM((to_integer(yCount - img_y) mod img_size_y),(to_integer(xCount - img_x)) mod img_size_x) when is_img_painted = '1' else (others => '0');
--    img_clr <= COLOR_GIF_ROM(to_integer(current_frame_gif(11 downto 6)), (to_integer(yCount - img_y) mod img_size_y),(to_integer(xCount - img_x)) mod img_size_x) when is_img_painted = '1' else (others => '0');
    img_clr <= apple_GIF_ROM(to_integer(current_frame_gif(11 downto 3)), (to_integer(yCount - img_y) mod 16),(to_integer(xCount - img_x)) mod 16) when is_img_painted = '1' else (others => '0');

    brick_clr <= BRICK_ROM((to_integer(yCount) mod 16),(to_integer(xCount) mod 16)) when border = '1' else (others => '0');

	snake_clr <= SNAKE_ROM((to_integer(yCount) mod 8),(to_integer(xCount) mod 8)) when snakeBody /= (127 downto 0 => '0') else (others => '0');

    vga_controller : entity work.vga_controller_640_60(Behavioral)
        Port map (rst => '0', pixel_clk => pixel_clk, HS => hsync, VS => vsync, hcount => xCount, vcount => yCount, blank => display);

    clk_div_unit_25Mhz : entity work.nbit_clk_div(Behavioral)
        Generic map (div_factor => 4,
                     high_count => 2,
                     num_of_bits => 3)
        Port map (clk_in => clk_100mhz, output => pixel_clk);

    -- instatiate random grid
    random_grid : entity work.randomGrid(Behavioral)
        Port map (pixel_clk => pixel_clk, rand_X => rand_X, rand_Y => rand_Y);

    update_clk : entity work.updateClk(Behavioral)
        Generic map (max_value => 4000000)
        Port map (clk_100mhz => clk_100mhz, update => update);

    up_sig : entity work.Debounce(Behavioral)
        Port map (clk => pixel_clk, rst => '0', noisy => btn_up, button_debounced => up);

    down_sig : entity work.Debounce(Behavioral)
        Port map (clk => pixel_clk, rst => '0', noisy => btn_down, button_debounced => down);

    left_sig : entity work.Debounce(Behavioral)
        Port map (clk => pixel_clk, rst => '0', noisy => btn_left, button_debounced => left);

    right_sig : entity work.Debounce(Behavioral)
        Port map (clk => pixel_clk, rst => '0', noisy => btn_right, button_debounced => right);

    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
        if pixel_clk = '1' then
            if start = '0' then
                snakeX(0) <= to_unsigned(40, 7);
                snakeY(0) <= to_unsigned(30, 7);
                for count in 1 to 127 loop
                    snakeX(count) <= to_unsigned(127, 7);
                    snakeY(count) <= to_unsigned(127, 7);
                end loop;
                size <= to_unsigned(1, 7);
                game_over <= '0';
            elsif game_over = '0' then
                if update = '1' then
                    for count in 1 to 127 loop
                        if size > count then
                            snakeX(count) <= snakeX(count-1);
                            snakeY(count) <= snakeY(count-1);
                        end if;
                    end loop;
                    case direction is
                        when "0001" =>
                            snakeY(0) <= snakeY(0) - to_unsigned(1, 7);
                        when "0010" =>
                            snakeY(0) <= snakeY(0) + to_unsigned(1, 7);
                        when "0100" =>
                            snakeX(0) <= snakeX(0) - to_unsigned(1, 7);
                        when "1000" =>
                            snakeX(0) <= snakeX(0) + to_unsigned(1, 7);
                        when others =>
                            null;
                    end case;
                else 
                    if img_clr /= "000000000000" and (snakeBody /= (127 downto 0 => '0')) then                    
--                    if (snakeX(0) = pearX) and (snakeY(0) = pearY) then
                        img_x <= rand_X & "0000";
                        img_y <= rand_Y & "0000";
                        if size < (128 - SIZE_INCREMENT) then
                            size <= size + SIZE_INCREMENT;
                        end if;
                    
                    -- elsif border = '1' and snakeBody(0) = '1' then
                    elsif brick_clr /= "000000000000" and snakeBody(0) = '1' then
                         game_over <= '1';
                    
                    elsif (snakeBody(127 downto 1) /= (127 downto 1 => '0') and snakeBody(0) = '1') then
                        game_over <= '1';
                    end if;
                end if;
            end if;
        end if;
        end if;
    end process;

    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
            if pixel_clk = '1' then
            if (up = '1' and direction /= "0010") then
                direction <= "0001";
            elsif (down = '1' and direction /= "0001") then
                direction <= "0010";
            elsif (left = '1' and  direction /= "1000") then
                direction <= "0100";
            elsif (right  = '1' and direction /= "0100") then
                direction <= "1000";
            end if;
            end if;
        end if;
    end process;

    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
        if pixel_clk = '1' then
            if switch(0) = '1' then
                if ((xCount(9 downto 3) = 0) or (xCount(9 downto 3) = 79) or (yCount(9 downto 3) = 0) or (yCount(9 downto 3) = 59) or ((xCount(9 downto 3) = 10) and (yCount(9 downto 3) >= 10 and yCount(9 downto 3) <= 20)) or ((xCount(9 downto 3) = 69) and (yCount(9 downto 3) >= 39 and yCount(9 downto 3) <= 49)) or ((yCount(9 downto 3) = 10) and (xCount(9 downto 3) >= 10 and xCount(9 downto 3) <= 20)) or ((yCount(9 downto 3) = 49) and (xCount(9 downto 3) >= 59 and xCount(9 downto 3) <= 69))) then
                    border <= '1';
                else 
                    border <= '0';
                end if;
            elsif switch(1) = '1' then
                if ((xCount(9 downto 3) = 0) or (xCount(9 downto 3) = 79) or (yCount(9 downto 3) = 0) or (yCount(9 downto 3) = 59) or((yCount(9 downto 3) = 20) and (xCount(9 downto 3) >= 10 and xCount(9 downto 3) <= 69)) or ((yCount(9 downto 3) =40 ) and (xCount(9 downto 3) >= 10 and xCount(9 downto 3) <= 69))) then
                    border <= '1';
                else 
                    border <= '0';
                end if;
            elsif switch(2) = '1' then
                if ((xCount(9 downto 3) = 0) or (xCount(9 downto 3) = 79) or (yCount(9 downto 3) = 0) or (yCount(9 downto 3) = 59) or ((xCount(9 downto 3) = 39) and (yCount(9 downto 3) >= 0 and yCount(9 downto 3) <=10)) or ((xCount(9 downto 3) = 39) and (yCount(9 downto 3) >= 49 and  yCount(9 downto 3)<=59))) then
                    border <= '1';
                else 
                    border <= '0';
                end if;
            else
                -- if (xCount(9 downto 3) = 0) or (xCount(9 downto 3) = 79) or (yCount(9 downto 3) = 0) or (yCount(9 downto 3) = 59) then
                if (xCount < img_size_x or xCount > 640 - img_size_x or yCount < img_size_y or yCount > 480 - img_size_y) then    
                    border <= '1';
                else 
                    border <= '0';
                end if;
            end if;
        end if;
        end if;
    end process;

    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
        if pixel_clk = '1' then
            if (xCount(9 downto 3) = pearX) and (yCount(9 downto 3) = pearY) then
                pear <= '1';
                
                
                -- pear <= ROM(to_integer(yCount(9 downto 3))) (to_integer(xCount(9 downto 3)));
            else
                pear <= '0';
            end if;
        end if;
        end if;
    end process;

    process(clk_100mhz)
    begin
        if rising_edge(clk_100mhz) then
        if pixel_clk = '1' then
            for count in 0 to 127 loop
                if (xCount(9 downto 3) = snakeX(count)) and (yCount(9 downto 3) = snakeY(count)) then
                    snakeBody(count) <= '1';
                else
                    snakeBody(count) <= '0';
                end if;
            end loop;
        end if;
        end if;
    end process;
    
    vgared <= rgb(11 downto 8);
    vgagreen <= rgb(7 downto 4);
    vgablue <= rgb(3 downto 0);
    
    rgb <= (others => '0') when display = '1' else 
           "111100000000" when game_over = '1' else
           snake_clr when (snakeBody /= (127 downto 0 => '0')) else
           brick_clr when border = '1' else 
           img_clr;

--    vgared <= "1111" when (display = '0' and (img_clr /= "000000000000" or game_over = '1')) else "0000";
--    vgagreen <= "1111" when display = '0' and (snakeBody /= (127 downto 0 => '0') and game_over = '0') ;
--    vgablue <= "1111" when (display = '0' and (border = '1' and game_over = '0')) else "0000";

end Behavioral;